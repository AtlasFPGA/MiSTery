
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"d9",x"c4",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c0",x"d9",x"c4"),
    14 => (x"48",x"f8",x"fe",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fc",x"f1"),
    19 => (x"fc",x"1e",x"87",x"fd"),
    20 => (x"ff",x"4a",x"71",x"86"),
    21 => (x"48",x"69",x"49",x"c0"),
    22 => (x"70",x"98",x"c0",x"c4"),
    23 => (x"02",x"98",x"48",x"7e"),
    24 => (x"79",x"72",x"87",x"f4"),
    25 => (x"26",x"8e",x"fc",x"48"),
    26 => (x"1e",x"72",x"1e",x"4f"),
    27 => (x"48",x"12",x"1e",x"73"),
    28 => (x"87",x"ca",x"02",x"11"),
    29 => (x"98",x"df",x"c3",x"4b"),
    30 => (x"02",x"88",x"73",x"9b"),
    31 => (x"4b",x"26",x"87",x"f0"),
    32 => (x"4f",x"26",x"4a",x"26"),
    33 => (x"72",x"1e",x"73",x"1e"),
    34 => (x"04",x"8b",x"c1",x"1e"),
    35 => (x"48",x"12",x"87",x"ca"),
    36 => (x"87",x"c4",x"02",x"11"),
    37 => (x"87",x"f1",x"02",x"88"),
    38 => (x"4b",x"26",x"4a",x"26"),
    39 => (x"74",x"1e",x"4f",x"26"),
    40 => (x"72",x"1e",x"73",x"1e"),
    41 => (x"04",x"8b",x"c1",x"1e"),
    42 => (x"48",x"12",x"87",x"d0"),
    43 => (x"87",x"ca",x"02",x"11"),
    44 => (x"98",x"df",x"c3",x"4c"),
    45 => (x"02",x"88",x"74",x"9c"),
    46 => (x"4a",x"26",x"87",x"eb"),
    47 => (x"4c",x"26",x"4b",x"26"),
    48 => (x"73",x"1e",x"4f",x"26"),
    49 => (x"a9",x"73",x"81",x"48"),
    50 => (x"12",x"87",x"c5",x"02"),
    51 => (x"87",x"f6",x"05",x"53"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"a9",x"73",x"81",x"48"),
    54 => (x"f9",x"53",x"72",x"05"),
    55 => (x"1e",x"4f",x"26",x"87"),
    56 => (x"9a",x"72",x"1e",x"73"),
    57 => (x"87",x"e7",x"c0",x"02"),
    58 => (x"4b",x"c1",x"48",x"c0"),
    59 => (x"d1",x"06",x"a9",x"72"),
    60 => (x"06",x"82",x"72",x"87"),
    61 => (x"83",x"73",x"87",x"c9"),
    62 => (x"f4",x"01",x"a9",x"72"),
    63 => (x"c1",x"87",x"c3",x"87"),
    64 => (x"a9",x"72",x"3a",x"b2"),
    65 => (x"80",x"73",x"89",x"03"),
    66 => (x"2b",x"2a",x"c1",x"07"),
    67 => (x"26",x"87",x"f3",x"05"),
    68 => (x"1e",x"4f",x"26",x"4b"),
    69 => (x"4d",x"c4",x"1e",x"75"),
    70 => (x"04",x"a1",x"b7",x"71"),
    71 => (x"81",x"c1",x"b9",x"ff"),
    72 => (x"72",x"07",x"bd",x"c3"),
    73 => (x"ff",x"04",x"a2",x"b7"),
    74 => (x"c1",x"82",x"c1",x"ba"),
    75 => (x"ee",x"fe",x"07",x"bd"),
    76 => (x"04",x"2d",x"c1",x"87"),
    77 => (x"80",x"c1",x"b8",x"ff"),
    78 => (x"ff",x"04",x"2d",x"07"),
    79 => (x"07",x"81",x"c1",x"b9"),
    80 => (x"4f",x"26",x"4d",x"26"),
    81 => (x"71",x"1e",x"73",x"1e"),
    82 => (x"4b",x"66",x"c8",x"4a"),
    83 => (x"71",x"8b",x"c1",x"49"),
    84 => (x"87",x"cf",x"02",x"99"),
    85 => (x"d4",x"ff",x"48",x"12"),
    86 => (x"49",x"73",x"78",x"08"),
    87 => (x"99",x"71",x"8b",x"c1"),
    88 => (x"26",x"87",x"f1",x"05"),
    89 => (x"0e",x"4f",x"26",x"4b"),
    90 => (x"0e",x"5c",x"5b",x"5e"),
    91 => (x"d4",x"ff",x"4a",x"71"),
    92 => (x"4b",x"66",x"cc",x"4c"),
    93 => (x"71",x"8b",x"c1",x"49"),
    94 => (x"87",x"ce",x"02",x"99"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"c1",x"49",x"73",x"52"),
    97 => (x"05",x"99",x"71",x"8b"),
    98 => (x"4c",x"26",x"87",x"f2"),
    99 => (x"4f",x"26",x"4b",x"26"),
   100 => (x"ff",x"1e",x"73",x"1e"),
   101 => (x"ff",x"c3",x"4b",x"d4"),
   102 => (x"c3",x"4a",x"6b",x"7b"),
   103 => (x"49",x"6b",x"7b",x"ff"),
   104 => (x"b1",x"72",x"32",x"c8"),
   105 => (x"6b",x"7b",x"ff",x"c3"),
   106 => (x"71",x"31",x"c8",x"4a"),
   107 => (x"7b",x"ff",x"c3",x"b2"),
   108 => (x"32",x"c8",x"49",x"6b"),
   109 => (x"48",x"71",x"b1",x"72"),
   110 => (x"4f",x"26",x"4b",x"26"),
   111 => (x"5c",x"5b",x"5e",x"0e"),
   112 => (x"4d",x"71",x"0e",x"5d"),
   113 => (x"75",x"4c",x"d4",x"ff"),
   114 => (x"98",x"ff",x"c3",x"48"),
   115 => (x"fe",x"c3",x"7c",x"70"),
   116 => (x"c8",x"05",x"bf",x"f8"),
   117 => (x"48",x"66",x"d0",x"87"),
   118 => (x"a6",x"d4",x"30",x"c9"),
   119 => (x"49",x"66",x"d0",x"58"),
   120 => (x"48",x"71",x"29",x"d8"),
   121 => (x"70",x"98",x"ff",x"c3"),
   122 => (x"49",x"66",x"d0",x"7c"),
   123 => (x"48",x"71",x"29",x"d0"),
   124 => (x"70",x"98",x"ff",x"c3"),
   125 => (x"49",x"66",x"d0",x"7c"),
   126 => (x"48",x"71",x"29",x"c8"),
   127 => (x"70",x"98",x"ff",x"c3"),
   128 => (x"48",x"66",x"d0",x"7c"),
   129 => (x"70",x"98",x"ff",x"c3"),
   130 => (x"d0",x"49",x"75",x"7c"),
   131 => (x"c3",x"48",x"71",x"29"),
   132 => (x"7c",x"70",x"98",x"ff"),
   133 => (x"f0",x"c9",x"4b",x"6c"),
   134 => (x"ff",x"c3",x"4a",x"ff"),
   135 => (x"87",x"cf",x"05",x"ab"),
   136 => (x"6c",x"7c",x"71",x"49"),
   137 => (x"02",x"8a",x"c1",x"4b"),
   138 => (x"ab",x"71",x"87",x"c5"),
   139 => (x"73",x"87",x"f2",x"02"),
   140 => (x"26",x"4d",x"26",x"48"),
   141 => (x"26",x"4b",x"26",x"4c"),
   142 => (x"49",x"c0",x"1e",x"4f"),
   143 => (x"c3",x"48",x"d4",x"ff"),
   144 => (x"81",x"c1",x"78",x"ff"),
   145 => (x"a9",x"b7",x"c8",x"c3"),
   146 => (x"26",x"87",x"f1",x"04"),
   147 => (x"5b",x"5e",x"0e",x"4f"),
   148 => (x"c0",x"0e",x"5d",x"5c"),
   149 => (x"f7",x"c1",x"f0",x"ff"),
   150 => (x"c0",x"c0",x"c1",x"4d"),
   151 => (x"4b",x"c0",x"c0",x"c0"),
   152 => (x"c4",x"87",x"d6",x"ff"),
   153 => (x"c0",x"4c",x"df",x"f8"),
   154 => (x"fd",x"49",x"75",x"1e"),
   155 => (x"86",x"c4",x"87",x"ce"),
   156 => (x"c0",x"05",x"a8",x"c1"),
   157 => (x"d4",x"ff",x"87",x"e5"),
   158 => (x"78",x"ff",x"c3",x"48"),
   159 => (x"e1",x"c0",x"1e",x"73"),
   160 => (x"49",x"e9",x"c1",x"f0"),
   161 => (x"c4",x"87",x"f5",x"fc"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"d4",x"ff",x"87",x"ca"),
   164 => (x"78",x"ff",x"c3",x"48"),
   165 => (x"87",x"cb",x"48",x"c1"),
   166 => (x"c1",x"87",x"de",x"fe"),
   167 => (x"c6",x"ff",x"05",x"8c"),
   168 => (x"26",x"48",x"c0",x"87"),
   169 => (x"26",x"4c",x"26",x"4d"),
   170 => (x"0e",x"4f",x"26",x"4b"),
   171 => (x"0e",x"5c",x"5b",x"5e"),
   172 => (x"c1",x"f0",x"ff",x"c0"),
   173 => (x"d4",x"ff",x"4c",x"c1"),
   174 => (x"78",x"ff",x"c3",x"48"),
   175 => (x"1e",x"c0",x"4b",x"d3"),
   176 => (x"f7",x"fb",x"49",x"74"),
   177 => (x"70",x"86",x"c4",x"87"),
   178 => (x"87",x"ca",x"05",x"98"),
   179 => (x"c3",x"48",x"d4",x"ff"),
   180 => (x"48",x"c1",x"78",x"ff"),
   181 => (x"e0",x"fd",x"87",x"ca"),
   182 => (x"05",x"8b",x"c1",x"87"),
   183 => (x"48",x"c0",x"87",x"e0"),
   184 => (x"4b",x"26",x"4c",x"26"),
   185 => (x"5e",x"0e",x"4f",x"26"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"c4",x"fd",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"fb",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"e0",x"fe"),
   195 => (x"87",x"e2",x"c1",x"48"),
   196 => (x"70",x"87",x"fd",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fe",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"c9"),
   201 => (x"75",x"87",x"cb",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"de",x"fc"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"fc",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"d5",x"48",x"c1",x"87"),
   215 => (x"d1",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"48",x"c0",x"87",x"c4"),
   218 => (x"8c",x"c1",x"87",x"c8"),
   219 => (x"87",x"fc",x"fe",x"05"),
   220 => (x"4d",x"26",x"48",x"c0"),
   221 => (x"4b",x"26",x"4c",x"26"),
   222 => (x"5e",x"0e",x"4f",x"26"),
   223 => (x"0e",x"5d",x"5c",x"5b"),
   224 => (x"c0",x"4d",x"d0",x"ff"),
   225 => (x"c0",x"c1",x"d0",x"e5"),
   226 => (x"f8",x"fe",x"c3",x"4c"),
   227 => (x"c7",x"78",x"c1",x"48"),
   228 => (x"fa",x"7d",x"c2",x"4b"),
   229 => (x"7d",x"c3",x"87",x"e3"),
   230 => (x"49",x"74",x"1e",x"c0"),
   231 => (x"c4",x"87",x"dd",x"f8"),
   232 => (x"05",x"a8",x"c1",x"86"),
   233 => (x"c2",x"4b",x"87",x"c1"),
   234 => (x"87",x"c5",x"05",x"ab"),
   235 => (x"f6",x"c0",x"48",x"c0"),
   236 => (x"05",x"8b",x"c1",x"87"),
   237 => (x"fc",x"87",x"da",x"ff"),
   238 => (x"fe",x"c3",x"87",x"ec"),
   239 => (x"98",x"70",x"58",x"fc"),
   240 => (x"c1",x"87",x"cd",x"05"),
   241 => (x"f0",x"ff",x"c0",x"1e"),
   242 => (x"f7",x"49",x"d0",x"c1"),
   243 => (x"86",x"c4",x"87",x"ee"),
   244 => (x"c3",x"48",x"d4",x"ff"),
   245 => (x"e8",x"c4",x"78",x"ff"),
   246 => (x"c0",x"ff",x"c3",x"87"),
   247 => (x"ff",x"7d",x"c2",x"58"),
   248 => (x"ff",x"c3",x"48",x"d4"),
   249 => (x"26",x"48",x"c1",x"78"),
   250 => (x"26",x"4c",x"26",x"4d"),
   251 => (x"0e",x"4f",x"26",x"4b"),
   252 => (x"5d",x"5c",x"5b",x"5e"),
   253 => (x"c3",x"4d",x"71",x"0e"),
   254 => (x"d4",x"ff",x"4c",x"ff"),
   255 => (x"ff",x"7b",x"74",x"4b"),
   256 => (x"c3",x"c4",x"48",x"d0"),
   257 => (x"75",x"7b",x"74",x"78"),
   258 => (x"f0",x"ff",x"c0",x"1e"),
   259 => (x"f6",x"49",x"d8",x"c1"),
   260 => (x"86",x"c4",x"87",x"ea"),
   261 => (x"c5",x"02",x"98",x"70"),
   262 => (x"c0",x"48",x"c1",x"87"),
   263 => (x"7b",x"74",x"87",x"ee"),
   264 => (x"c8",x"7b",x"fe",x"c3"),
   265 => (x"66",x"d4",x"1e",x"c0"),
   266 => (x"87",x"d8",x"f4",x"49"),
   267 => (x"7b",x"74",x"86",x"c4"),
   268 => (x"7b",x"74",x"7b",x"74"),
   269 => (x"4a",x"e0",x"da",x"d8"),
   270 => (x"05",x"6b",x"7b",x"74"),
   271 => (x"8a",x"c1",x"87",x"c5"),
   272 => (x"74",x"87",x"f5",x"05"),
   273 => (x"48",x"d0",x"ff",x"7b"),
   274 => (x"48",x"c0",x"78",x"c2"),
   275 => (x"4c",x"26",x"4d",x"26"),
   276 => (x"4f",x"26",x"4b",x"26"),
   277 => (x"5c",x"5b",x"5e",x"0e"),
   278 => (x"86",x"fc",x"0e",x"5d"),
   279 => (x"d4",x"ff",x"4b",x"71"),
   280 => (x"c5",x"7e",x"c0",x"4c"),
   281 => (x"4a",x"df",x"cd",x"ee"),
   282 => (x"6c",x"7c",x"ff",x"c3"),
   283 => (x"a8",x"fe",x"c3",x"48"),
   284 => (x"87",x"f8",x"c0",x"05"),
   285 => (x"9b",x"73",x"4d",x"74"),
   286 => (x"d4",x"87",x"cc",x"02"),
   287 => (x"49",x"73",x"1e",x"66"),
   288 => (x"c4",x"87",x"e4",x"f3"),
   289 => (x"ff",x"87",x"d4",x"86"),
   290 => (x"d1",x"c4",x"48",x"d0"),
   291 => (x"4a",x"66",x"d4",x"78"),
   292 => (x"c1",x"7d",x"ff",x"c3"),
   293 => (x"87",x"f8",x"05",x"8a"),
   294 => (x"c3",x"5a",x"a6",x"d8"),
   295 => (x"73",x"7c",x"7c",x"ff"),
   296 => (x"87",x"c5",x"05",x"9b"),
   297 => (x"d0",x"48",x"d0",x"ff"),
   298 => (x"7e",x"4a",x"c1",x"78"),
   299 => (x"fe",x"05",x"8a",x"c1"),
   300 => (x"48",x"6e",x"87",x"f6"),
   301 => (x"4d",x"26",x"8e",x"fc"),
   302 => (x"4b",x"26",x"4c",x"26"),
   303 => (x"73",x"1e",x"4f",x"26"),
   304 => (x"c0",x"4a",x"71",x"1e"),
   305 => (x"48",x"d4",x"ff",x"4b"),
   306 => (x"ff",x"78",x"ff",x"c3"),
   307 => (x"c3",x"c4",x"48",x"d0"),
   308 => (x"48",x"d4",x"ff",x"78"),
   309 => (x"72",x"78",x"ff",x"c3"),
   310 => (x"f0",x"ff",x"c0",x"1e"),
   311 => (x"f3",x"49",x"d1",x"c1"),
   312 => (x"86",x"c4",x"87",x"da"),
   313 => (x"d2",x"05",x"98",x"70"),
   314 => (x"1e",x"c0",x"c8",x"87"),
   315 => (x"fd",x"49",x"66",x"cc"),
   316 => (x"86",x"c4",x"87",x"e2"),
   317 => (x"d0",x"ff",x"4b",x"70"),
   318 => (x"73",x"78",x"c2",x"48"),
   319 => (x"26",x"4b",x"26",x"48"),
   320 => (x"5b",x"5e",x"0e",x"4f"),
   321 => (x"c0",x"0e",x"5d",x"5c"),
   322 => (x"f0",x"ff",x"c0",x"1e"),
   323 => (x"f2",x"49",x"c9",x"c1"),
   324 => (x"1e",x"d2",x"87",x"ea"),
   325 => (x"49",x"c0",x"ff",x"c3"),
   326 => (x"c8",x"87",x"f9",x"fc"),
   327 => (x"c1",x"4c",x"c0",x"86"),
   328 => (x"ac",x"b7",x"d2",x"84"),
   329 => (x"c3",x"87",x"f8",x"04"),
   330 => (x"bf",x"97",x"c0",x"ff"),
   331 => (x"99",x"c0",x"c3",x"49"),
   332 => (x"05",x"a9",x"c0",x"c1"),
   333 => (x"c3",x"87",x"e7",x"c0"),
   334 => (x"bf",x"97",x"c7",x"ff"),
   335 => (x"c3",x"31",x"d0",x"49"),
   336 => (x"bf",x"97",x"c8",x"ff"),
   337 => (x"72",x"32",x"c8",x"4a"),
   338 => (x"c9",x"ff",x"c3",x"b1"),
   339 => (x"b1",x"4a",x"bf",x"97"),
   340 => (x"ff",x"cf",x"4c",x"71"),
   341 => (x"c1",x"9c",x"ff",x"ff"),
   342 => (x"c1",x"34",x"ca",x"84"),
   343 => (x"ff",x"c3",x"87",x"e7"),
   344 => (x"49",x"bf",x"97",x"c9"),
   345 => (x"99",x"c6",x"31",x"c1"),
   346 => (x"97",x"ca",x"ff",x"c3"),
   347 => (x"b7",x"c7",x"4a",x"bf"),
   348 => (x"c3",x"b1",x"72",x"2a"),
   349 => (x"bf",x"97",x"c5",x"ff"),
   350 => (x"9d",x"cf",x"4d",x"4a"),
   351 => (x"97",x"c6",x"ff",x"c3"),
   352 => (x"9a",x"c3",x"4a",x"bf"),
   353 => (x"ff",x"c3",x"32",x"ca"),
   354 => (x"4b",x"bf",x"97",x"c7"),
   355 => (x"b2",x"73",x"33",x"c2"),
   356 => (x"97",x"c8",x"ff",x"c3"),
   357 => (x"c0",x"c3",x"4b",x"bf"),
   358 => (x"2b",x"b7",x"c6",x"9b"),
   359 => (x"81",x"c2",x"b2",x"73"),
   360 => (x"30",x"71",x"48",x"c1"),
   361 => (x"48",x"c1",x"49",x"70"),
   362 => (x"4d",x"70",x"30",x"75"),
   363 => (x"84",x"c1",x"4c",x"72"),
   364 => (x"c0",x"c8",x"94",x"71"),
   365 => (x"cc",x"06",x"ad",x"b7"),
   366 => (x"b7",x"34",x"c1",x"87"),
   367 => (x"b7",x"c0",x"c8",x"2d"),
   368 => (x"f4",x"ff",x"01",x"ad"),
   369 => (x"26",x"48",x"74",x"87"),
   370 => (x"26",x"4c",x"26",x"4d"),
   371 => (x"0e",x"4f",x"26",x"4b"),
   372 => (x"5d",x"5c",x"5b",x"5e"),
   373 => (x"c4",x"86",x"f8",x"0e"),
   374 => (x"c0",x"48",x"e8",x"c7"),
   375 => (x"e0",x"ff",x"c3",x"78"),
   376 => (x"fb",x"49",x"c0",x"1e"),
   377 => (x"86",x"c4",x"87",x"d8"),
   378 => (x"c5",x"05",x"98",x"70"),
   379 => (x"c9",x"48",x"c0",x"87"),
   380 => (x"4d",x"c0",x"87",x"c0"),
   381 => (x"c2",x"c1",x"7e",x"c1"),
   382 => (x"c4",x"49",x"bf",x"d4"),
   383 => (x"71",x"4a",x"d6",x"c0"),
   384 => (x"ff",x"e9",x"4b",x"c8"),
   385 => (x"05",x"98",x"70",x"87"),
   386 => (x"7e",x"c0",x"87",x"c2"),
   387 => (x"bf",x"d0",x"c2",x"c1"),
   388 => (x"f2",x"c0",x"c4",x"49"),
   389 => (x"4b",x"c8",x"71",x"4a"),
   390 => (x"70",x"87",x"e9",x"e9"),
   391 => (x"87",x"c2",x"05",x"98"),
   392 => (x"02",x"6e",x"7e",x"c0"),
   393 => (x"c4",x"87",x"fd",x"c0"),
   394 => (x"4d",x"bf",x"e6",x"c6"),
   395 => (x"9f",x"de",x"c7",x"c4"),
   396 => (x"c5",x"48",x"7e",x"bf"),
   397 => (x"05",x"a8",x"ea",x"d6"),
   398 => (x"c6",x"c4",x"87",x"c7"),
   399 => (x"ce",x"4d",x"bf",x"e6"),
   400 => (x"ca",x"48",x"6e",x"87"),
   401 => (x"02",x"a8",x"d5",x"e9"),
   402 => (x"48",x"c0",x"87",x"c5"),
   403 => (x"c3",x"87",x"e3",x"c7"),
   404 => (x"75",x"1e",x"e0",x"ff"),
   405 => (x"87",x"e6",x"f9",x"49"),
   406 => (x"98",x"70",x"86",x"c4"),
   407 => (x"c0",x"87",x"c5",x"05"),
   408 => (x"87",x"ce",x"c7",x"48"),
   409 => (x"bf",x"d0",x"c2",x"c1"),
   410 => (x"f2",x"c0",x"c4",x"49"),
   411 => (x"4b",x"c8",x"71",x"4a"),
   412 => (x"70",x"87",x"d1",x"e8"),
   413 => (x"87",x"c8",x"05",x"98"),
   414 => (x"48",x"e8",x"c7",x"c4"),
   415 => (x"87",x"da",x"78",x"c1"),
   416 => (x"bf",x"d4",x"c2",x"c1"),
   417 => (x"d6",x"c0",x"c4",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"f5",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c6",x"48",x"c0",x"87"),
   422 => (x"c7",x"c4",x"87",x"d8"),
   423 => (x"49",x"bf",x"97",x"de"),
   424 => (x"05",x"a9",x"d5",x"c1"),
   425 => (x"c4",x"87",x"cd",x"c0"),
   426 => (x"bf",x"97",x"df",x"c7"),
   427 => (x"a9",x"ea",x"c2",x"49"),
   428 => (x"87",x"c5",x"c0",x"02"),
   429 => (x"f9",x"c5",x"48",x"c0"),
   430 => (x"e0",x"ff",x"c3",x"87"),
   431 => (x"48",x"7e",x"bf",x"97"),
   432 => (x"02",x"a8",x"e9",x"c3"),
   433 => (x"6e",x"87",x"ce",x"c0"),
   434 => (x"a8",x"eb",x"c3",x"48"),
   435 => (x"87",x"c5",x"c0",x"02"),
   436 => (x"dd",x"c5",x"48",x"c0"),
   437 => (x"eb",x"ff",x"c3",x"87"),
   438 => (x"99",x"49",x"bf",x"97"),
   439 => (x"87",x"cc",x"c0",x"05"),
   440 => (x"97",x"ec",x"ff",x"c3"),
   441 => (x"a9",x"c2",x"49",x"bf"),
   442 => (x"87",x"c5",x"c0",x"02"),
   443 => (x"c1",x"c5",x"48",x"c0"),
   444 => (x"ed",x"ff",x"c3",x"87"),
   445 => (x"c4",x"48",x"bf",x"97"),
   446 => (x"70",x"58",x"e4",x"c7"),
   447 => (x"88",x"c1",x"48",x"4c"),
   448 => (x"58",x"e8",x"c7",x"c4"),
   449 => (x"97",x"ee",x"ff",x"c3"),
   450 => (x"81",x"75",x"49",x"bf"),
   451 => (x"97",x"ef",x"ff",x"c3"),
   452 => (x"32",x"c8",x"4a",x"bf"),
   453 => (x"c4",x"7e",x"a1",x"72"),
   454 => (x"6e",x"48",x"f8",x"cb"),
   455 => (x"f0",x"ff",x"c3",x"78"),
   456 => (x"c8",x"48",x"bf",x"97"),
   457 => (x"c7",x"c4",x"58",x"a6"),
   458 => (x"c2",x"02",x"bf",x"e8"),
   459 => (x"c2",x"c1",x"87",x"cf"),
   460 => (x"c4",x"49",x"bf",x"d0"),
   461 => (x"71",x"4a",x"f2",x"c0"),
   462 => (x"c7",x"e5",x"4b",x"c8"),
   463 => (x"02",x"98",x"70",x"87"),
   464 => (x"c0",x"87",x"c5",x"c0"),
   465 => (x"87",x"ea",x"c3",x"48"),
   466 => (x"bf",x"e0",x"c7",x"c4"),
   467 => (x"cc",x"cc",x"c4",x"4c"),
   468 => (x"c5",x"c0",x"c4",x"5c"),
   469 => (x"c8",x"49",x"bf",x"97"),
   470 => (x"c4",x"c0",x"c4",x"31"),
   471 => (x"a1",x"4a",x"bf",x"97"),
   472 => (x"c6",x"c0",x"c4",x"49"),
   473 => (x"d0",x"4a",x"bf",x"97"),
   474 => (x"49",x"a1",x"72",x"32"),
   475 => (x"97",x"c7",x"c0",x"c4"),
   476 => (x"32",x"d8",x"4a",x"bf"),
   477 => (x"c4",x"49",x"a1",x"72"),
   478 => (x"cb",x"c4",x"91",x"66"),
   479 => (x"c4",x"81",x"bf",x"f8"),
   480 => (x"c4",x"59",x"c0",x"cc"),
   481 => (x"bf",x"97",x"cd",x"c0"),
   482 => (x"c4",x"32",x"c8",x"4a"),
   483 => (x"bf",x"97",x"cc",x"c0"),
   484 => (x"c4",x"4a",x"a2",x"4b"),
   485 => (x"bf",x"97",x"ce",x"c0"),
   486 => (x"73",x"33",x"d0",x"4b"),
   487 => (x"c0",x"c4",x"4a",x"a2"),
   488 => (x"4b",x"bf",x"97",x"cf"),
   489 => (x"33",x"d8",x"9b",x"cf"),
   490 => (x"c4",x"4a",x"a2",x"73"),
   491 => (x"c2",x"5a",x"c4",x"cc"),
   492 => (x"c4",x"92",x"74",x"8a"),
   493 => (x"72",x"48",x"c4",x"cc"),
   494 => (x"c1",x"c1",x"78",x"a1"),
   495 => (x"f2",x"ff",x"c3",x"87"),
   496 => (x"c8",x"49",x"bf",x"97"),
   497 => (x"f1",x"ff",x"c3",x"31"),
   498 => (x"a1",x"4a",x"bf",x"97"),
   499 => (x"c7",x"31",x"c5",x"49"),
   500 => (x"29",x"c9",x"81",x"ff"),
   501 => (x"59",x"cc",x"cc",x"c4"),
   502 => (x"97",x"f7",x"ff",x"c3"),
   503 => (x"32",x"c8",x"4a",x"bf"),
   504 => (x"97",x"f6",x"ff",x"c3"),
   505 => (x"4a",x"a2",x"4b",x"bf"),
   506 => (x"6e",x"92",x"66",x"c4"),
   507 => (x"c8",x"cc",x"c4",x"82"),
   508 => (x"c0",x"cc",x"c4",x"5a"),
   509 => (x"c4",x"78",x"c0",x"48"),
   510 => (x"72",x"48",x"fc",x"cb"),
   511 => (x"cc",x"c4",x"78",x"a1"),
   512 => (x"cc",x"c4",x"48",x"cc"),
   513 => (x"c4",x"78",x"bf",x"c0"),
   514 => (x"c4",x"48",x"d0",x"cc"),
   515 => (x"78",x"bf",x"c4",x"cc"),
   516 => (x"bf",x"e8",x"c7",x"c4"),
   517 => (x"87",x"c9",x"c0",x"02"),
   518 => (x"30",x"c4",x"48",x"74"),
   519 => (x"c9",x"c0",x"7e",x"70"),
   520 => (x"c8",x"cc",x"c4",x"87"),
   521 => (x"30",x"c4",x"48",x"bf"),
   522 => (x"c7",x"c4",x"7e",x"70"),
   523 => (x"78",x"6e",x"48",x"ec"),
   524 => (x"8e",x"f8",x"48",x"c1"),
   525 => (x"4c",x"26",x"4d",x"26"),
   526 => (x"4f",x"26",x"4b",x"26"),
   527 => (x"5c",x"5b",x"5e",x"0e"),
   528 => (x"4a",x"71",x"0e",x"5d"),
   529 => (x"bf",x"e8",x"c7",x"c4"),
   530 => (x"72",x"87",x"cb",x"02"),
   531 => (x"72",x"2b",x"c7",x"4b"),
   532 => (x"9d",x"ff",x"c1",x"4d"),
   533 => (x"4b",x"72",x"87",x"c9"),
   534 => (x"4d",x"72",x"2b",x"c8"),
   535 => (x"c4",x"9d",x"ff",x"c3"),
   536 => (x"83",x"bf",x"f8",x"cb"),
   537 => (x"bf",x"cc",x"c2",x"c1"),
   538 => (x"87",x"d9",x"02",x"ab"),
   539 => (x"5b",x"d0",x"c2",x"c1"),
   540 => (x"1e",x"e0",x"ff",x"c3"),
   541 => (x"c5",x"f1",x"49",x"73"),
   542 => (x"70",x"86",x"c4",x"87"),
   543 => (x"87",x"c5",x"05",x"98"),
   544 => (x"e6",x"c0",x"48",x"c0"),
   545 => (x"e8",x"c7",x"c4",x"87"),
   546 => (x"87",x"d2",x"02",x"bf"),
   547 => (x"91",x"c4",x"49",x"75"),
   548 => (x"81",x"e0",x"ff",x"c3"),
   549 => (x"ff",x"cf",x"4c",x"69"),
   550 => (x"9c",x"ff",x"ff",x"ff"),
   551 => (x"49",x"75",x"87",x"cb"),
   552 => (x"ff",x"c3",x"91",x"c2"),
   553 => (x"69",x"9f",x"81",x"e0"),
   554 => (x"26",x"48",x"74",x"4c"),
   555 => (x"26",x"4c",x"26",x"4d"),
   556 => (x"0e",x"4f",x"26",x"4b"),
   557 => (x"5d",x"5c",x"5b",x"5e"),
   558 => (x"cc",x"86",x"f0",x"0e"),
   559 => (x"66",x"c8",x"59",x"a6"),
   560 => (x"c0",x"87",x"c5",x"05"),
   561 => (x"87",x"c5",x"c4",x"48"),
   562 => (x"c8",x"48",x"66",x"c8"),
   563 => (x"48",x"7e",x"70",x"80"),
   564 => (x"e0",x"c0",x"78",x"c0"),
   565 => (x"87",x"c8",x"02",x"66"),
   566 => (x"97",x"66",x"e0",x"c0"),
   567 => (x"87",x"c5",x"05",x"bf"),
   568 => (x"e8",x"c3",x"48",x"c0"),
   569 => (x"c1",x"1e",x"c0",x"87"),
   570 => (x"c4",x"d1",x"49",x"49"),
   571 => (x"70",x"86",x"c4",x"87"),
   572 => (x"c0",x"02",x"9c",x"4c"),
   573 => (x"c7",x"c4",x"87",x"fe"),
   574 => (x"e0",x"c0",x"4a",x"f0"),
   575 => (x"dd",x"ff",x"49",x"66"),
   576 => (x"98",x"70",x"87",x"e7"),
   577 => (x"87",x"ec",x"c0",x"02"),
   578 => (x"e0",x"c0",x"4a",x"74"),
   579 => (x"4b",x"cb",x"49",x"66"),
   580 => (x"87",x"ca",x"de",x"ff"),
   581 => (x"db",x"02",x"98",x"70"),
   582 => (x"74",x"1e",x"c0",x"87"),
   583 => (x"87",x"c4",x"02",x"9c"),
   584 => (x"87",x"c2",x"4d",x"c0"),
   585 => (x"49",x"75",x"4d",x"c1"),
   586 => (x"c4",x"87",x"c6",x"d0"),
   587 => (x"9c",x"4c",x"70",x"86"),
   588 => (x"87",x"c2",x"ff",x"05"),
   589 => (x"c2",x"02",x"9c",x"74"),
   590 => (x"a4",x"dc",x"87",x"d1"),
   591 => (x"69",x"48",x"6e",x"49"),
   592 => (x"49",x"a4",x"da",x"78"),
   593 => (x"c4",x"48",x"66",x"c8"),
   594 => (x"58",x"a6",x"c8",x"80"),
   595 => (x"c4",x"48",x"69",x"9f"),
   596 => (x"c4",x"78",x"08",x"66"),
   597 => (x"02",x"bf",x"e8",x"c7"),
   598 => (x"a4",x"d4",x"87",x"d2"),
   599 => (x"49",x"69",x"9f",x"49"),
   600 => (x"99",x"ff",x"ff",x"c0"),
   601 => (x"30",x"d0",x"48",x"71"),
   602 => (x"87",x"c5",x"58",x"a6"),
   603 => (x"c0",x"48",x"a6",x"cc"),
   604 => (x"49",x"66",x"cc",x"78"),
   605 => (x"bf",x"66",x"c4",x"48"),
   606 => (x"08",x"66",x"c4",x"80"),
   607 => (x"48",x"66",x"c8",x"78"),
   608 => (x"66",x"c8",x"78",x"c0"),
   609 => (x"c4",x"81",x"cc",x"49"),
   610 => (x"c8",x"79",x"bf",x"66"),
   611 => (x"81",x"d0",x"49",x"66"),
   612 => (x"c4",x"4d",x"79",x"c0"),
   613 => (x"66",x"c8",x"4c",x"66"),
   614 => (x"75",x"82",x"d4",x"4a"),
   615 => (x"72",x"91",x"c8",x"49"),
   616 => (x"41",x"c0",x"49",x"a1"),
   617 => (x"85",x"c1",x"79",x"6c"),
   618 => (x"04",x"ad",x"b7",x"c6"),
   619 => (x"6e",x"87",x"e7",x"ff"),
   620 => (x"2a",x"c9",x"4a",x"bf"),
   621 => (x"f0",x"c0",x"49",x"72"),
   622 => (x"e2",x"dc",x"ff",x"4a"),
   623 => (x"c8",x"4a",x"70",x"87"),
   624 => (x"c4",x"c1",x"49",x"66"),
   625 => (x"c1",x"79",x"72",x"81"),
   626 => (x"c0",x"87",x"c2",x"48"),
   627 => (x"26",x"8e",x"f0",x"48"),
   628 => (x"26",x"4c",x"26",x"4d"),
   629 => (x"0e",x"4f",x"26",x"4b"),
   630 => (x"5d",x"5c",x"5b",x"5e"),
   631 => (x"9c",x"4c",x"71",x"0e"),
   632 => (x"87",x"cb",x"c1",x"02"),
   633 => (x"69",x"49",x"a4",x"c8"),
   634 => (x"87",x"c3",x"c1",x"02"),
   635 => (x"6c",x"4a",x"66",x"d0"),
   636 => (x"48",x"a6",x"d0",x"49"),
   637 => (x"4d",x"78",x"a1",x"72"),
   638 => (x"e4",x"c7",x"c4",x"b9"),
   639 => (x"ba",x"ff",x"4a",x"bf"),
   640 => (x"99",x"71",x"99",x"72"),
   641 => (x"87",x"e4",x"c0",x"02"),
   642 => (x"6b",x"4b",x"a4",x"c4"),
   643 => (x"87",x"ec",x"f8",x"49"),
   644 => (x"c7",x"c4",x"7b",x"70"),
   645 => (x"6c",x"49",x"bf",x"e0"),
   646 => (x"75",x"7c",x"71",x"81"),
   647 => (x"e4",x"c7",x"c4",x"b9"),
   648 => (x"ba",x"ff",x"4a",x"bf"),
   649 => (x"99",x"71",x"99",x"72"),
   650 => (x"87",x"dc",x"ff",x"05"),
   651 => (x"26",x"7c",x"66",x"d0"),
   652 => (x"26",x"4c",x"26",x"4d"),
   653 => (x"1e",x"4f",x"26",x"4b"),
   654 => (x"4b",x"71",x"1e",x"73"),
   655 => (x"87",x"c7",x"02",x"9b"),
   656 => (x"69",x"49",x"a3",x"c8"),
   657 => (x"c0",x"87",x"c5",x"05"),
   658 => (x"87",x"f6",x"c0",x"48"),
   659 => (x"bf",x"fc",x"cb",x"c4"),
   660 => (x"4a",x"a3",x"c4",x"49"),
   661 => (x"8a",x"c2",x"4a",x"6a"),
   662 => (x"bf",x"e0",x"c7",x"c4"),
   663 => (x"49",x"a1",x"72",x"92"),
   664 => (x"bf",x"e4",x"c7",x"c4"),
   665 => (x"72",x"9a",x"6b",x"4a"),
   666 => (x"c2",x"c1",x"49",x"a1"),
   667 => (x"66",x"c8",x"59",x"d0"),
   668 => (x"c9",x"e9",x"71",x"1e"),
   669 => (x"70",x"86",x"c4",x"87"),
   670 => (x"87",x"c4",x"05",x"98"),
   671 => (x"87",x"c2",x"48",x"c0"),
   672 => (x"4b",x"26",x"48",x"c1"),
   673 => (x"73",x"1e",x"4f",x"26"),
   674 => (x"9b",x"4b",x"71",x"1e"),
   675 => (x"c8",x"87",x"c7",x"02"),
   676 => (x"05",x"69",x"49",x"a3"),
   677 => (x"48",x"c0",x"87",x"c5"),
   678 => (x"c4",x"87",x"f6",x"c0"),
   679 => (x"49",x"bf",x"fc",x"cb"),
   680 => (x"6a",x"4a",x"a3",x"c4"),
   681 => (x"c4",x"8a",x"c2",x"4a"),
   682 => (x"92",x"bf",x"e0",x"c7"),
   683 => (x"c4",x"49",x"a1",x"72"),
   684 => (x"4a",x"bf",x"e4",x"c7"),
   685 => (x"a1",x"72",x"9a",x"6b"),
   686 => (x"d0",x"c2",x"c1",x"49"),
   687 => (x"1e",x"66",x"c8",x"59"),
   688 => (x"87",x"eb",x"e4",x"71"),
   689 => (x"98",x"70",x"86",x"c4"),
   690 => (x"c0",x"87",x"c4",x"05"),
   691 => (x"c1",x"87",x"c2",x"48"),
   692 => (x"26",x"4b",x"26",x"48"),
   693 => (x"5b",x"5e",x"0e",x"4f"),
   694 => (x"f8",x"0e",x"5d",x"5c"),
   695 => (x"c4",x"7e",x"71",x"86"),
   696 => (x"78",x"ff",x"48",x"a6"),
   697 => (x"ff",x"ff",x"ff",x"c1"),
   698 => (x"c0",x"4d",x"ff",x"ff"),
   699 => (x"d4",x"4a",x"6e",x"4b"),
   700 => (x"c8",x"49",x"73",x"82"),
   701 => (x"49",x"a1",x"72",x"91"),
   702 => (x"69",x"4c",x"66",x"d8"),
   703 => (x"ac",x"b7",x"c0",x"8c"),
   704 => (x"75",x"87",x"cb",x"04"),
   705 => (x"c5",x"03",x"ac",x"b7"),
   706 => (x"5b",x"a6",x"c8",x"87"),
   707 => (x"83",x"c1",x"4d",x"74"),
   708 => (x"04",x"ab",x"b7",x"c6"),
   709 => (x"c4",x"87",x"d6",x"ff"),
   710 => (x"8e",x"f8",x"48",x"66"),
   711 => (x"4c",x"26",x"4d",x"26"),
   712 => (x"4f",x"26",x"4b",x"26"),
   713 => (x"5c",x"5b",x"5e",x"0e"),
   714 => (x"86",x"f0",x"0e",x"5d"),
   715 => (x"a6",x"c4",x"7e",x"71"),
   716 => (x"ff",x"ff",x"c1",x"48"),
   717 => (x"78",x"ff",x"ff",x"ff"),
   718 => (x"78",x"ff",x"80",x"c4"),
   719 => (x"4c",x"c0",x"4d",x"c0"),
   720 => (x"83",x"d4",x"4b",x"6e"),
   721 => (x"92",x"c8",x"4a",x"74"),
   722 => (x"75",x"4a",x"a2",x"73"),
   723 => (x"73",x"91",x"c8",x"49"),
   724 => (x"48",x"6a",x"49",x"a1"),
   725 => (x"a6",x"d0",x"88",x"69"),
   726 => (x"02",x"ad",x"74",x"58"),
   727 => (x"66",x"c4",x"87",x"cf"),
   728 => (x"87",x"c9",x"03",x"a8"),
   729 => (x"c4",x"5c",x"a6",x"cc"),
   730 => (x"66",x"cc",x"48",x"a6"),
   731 => (x"c6",x"84",x"c1",x"78"),
   732 => (x"ff",x"04",x"ac",x"b7"),
   733 => (x"85",x"c1",x"87",x"ca"),
   734 => (x"04",x"ad",x"b7",x"c6"),
   735 => (x"c8",x"87",x"ff",x"fe"),
   736 => (x"8e",x"f0",x"48",x"66"),
   737 => (x"4c",x"26",x"4d",x"26"),
   738 => (x"4f",x"26",x"4b",x"26"),
   739 => (x"5c",x"5b",x"5e",x"0e"),
   740 => (x"86",x"ec",x"0e",x"5d"),
   741 => (x"e4",x"c0",x"4b",x"71"),
   742 => (x"28",x"c9",x"48",x"66"),
   743 => (x"c4",x"58",x"a6",x"c8"),
   744 => (x"4a",x"bf",x"e4",x"c7"),
   745 => (x"48",x"72",x"ba",x"ff"),
   746 => (x"cc",x"98",x"66",x"c4"),
   747 => (x"9b",x"73",x"58",x"a6"),
   748 => (x"87",x"c1",x"c3",x"02"),
   749 => (x"69",x"49",x"a3",x"c8"),
   750 => (x"87",x"f9",x"c2",x"02"),
   751 => (x"98",x"6b",x"48",x"72"),
   752 => (x"c4",x"58",x"a6",x"d4"),
   753 => (x"7e",x"6c",x"4c",x"a3"),
   754 => (x"d0",x"48",x"66",x"c8"),
   755 => (x"c6",x"05",x"a8",x"66"),
   756 => (x"7b",x"66",x"c4",x"87"),
   757 => (x"c8",x"87",x"cc",x"c2"),
   758 => (x"49",x"73",x"1e",x"66"),
   759 => (x"c4",x"87",x"f6",x"fb"),
   760 => (x"c0",x"4d",x"70",x"86"),
   761 => (x"d0",x"04",x"ad",x"b7"),
   762 => (x"4a",x"a3",x"d4",x"87"),
   763 => (x"91",x"c8",x"49",x"75"),
   764 => (x"21",x"49",x"a1",x"72"),
   765 => (x"c7",x"7c",x"69",x"7b"),
   766 => (x"cc",x"7b",x"c0",x"87"),
   767 => (x"7c",x"69",x"49",x"a3"),
   768 => (x"6b",x"48",x"66",x"c4"),
   769 => (x"58",x"a6",x"c8",x"88"),
   770 => (x"73",x"1e",x"66",x"d0"),
   771 => (x"87",x"c5",x"fb",x"49"),
   772 => (x"4d",x"70",x"86",x"c4"),
   773 => (x"49",x"a3",x"c4",x"c1"),
   774 => (x"69",x"48",x"a6",x"c8"),
   775 => (x"48",x"66",x"d0",x"78"),
   776 => (x"06",x"a8",x"66",x"c8"),
   777 => (x"c0",x"87",x"f2",x"c0"),
   778 => (x"c0",x"04",x"ad",x"b7"),
   779 => (x"a6",x"cc",x"87",x"eb"),
   780 => (x"78",x"a3",x"d4",x"48"),
   781 => (x"91",x"c8",x"49",x"75"),
   782 => (x"d0",x"81",x"66",x"cc"),
   783 => (x"88",x"69",x"48",x"66"),
   784 => (x"66",x"c8",x"49",x"70"),
   785 => (x"87",x"d1",x"06",x"a9"),
   786 => (x"d7",x"fb",x"49",x"73"),
   787 => (x"c8",x"49",x"70",x"87"),
   788 => (x"81",x"66",x"cc",x"91"),
   789 => (x"6e",x"41",x"66",x"d0"),
   790 => (x"1e",x"66",x"c4",x"79"),
   791 => (x"f6",x"f5",x"49",x"73"),
   792 => (x"c3",x"86",x"c4",x"87"),
   793 => (x"73",x"1e",x"e0",x"ff"),
   794 => (x"87",x"cb",x"f7",x"49"),
   795 => (x"a3",x"d0",x"86",x"c4"),
   796 => (x"66",x"e4",x"c0",x"49"),
   797 => (x"26",x"8e",x"ec",x"79"),
   798 => (x"26",x"4c",x"26",x"4d"),
   799 => (x"1e",x"4f",x"26",x"4b"),
   800 => (x"4b",x"71",x"1e",x"73"),
   801 => (x"e4",x"c0",x"02",x"9b"),
   802 => (x"d0",x"cc",x"c4",x"87"),
   803 => (x"c2",x"4a",x"73",x"5b"),
   804 => (x"e0",x"c7",x"c4",x"8a"),
   805 => (x"c4",x"92",x"49",x"bf"),
   806 => (x"48",x"bf",x"fc",x"cb"),
   807 => (x"cc",x"c4",x"80",x"72"),
   808 => (x"48",x"71",x"58",x"d4"),
   809 => (x"c7",x"c4",x"30",x"c4"),
   810 => (x"ed",x"c0",x"58",x"f0"),
   811 => (x"cc",x"cc",x"c4",x"87"),
   812 => (x"c0",x"cc",x"c4",x"48"),
   813 => (x"cc",x"c4",x"78",x"bf"),
   814 => (x"cc",x"c4",x"48",x"d0"),
   815 => (x"c4",x"78",x"bf",x"c4"),
   816 => (x"02",x"bf",x"e8",x"c7"),
   817 => (x"c7",x"c4",x"87",x"c9"),
   818 => (x"c4",x"49",x"bf",x"e0"),
   819 => (x"c4",x"87",x"c7",x"31"),
   820 => (x"49",x"bf",x"c8",x"cc"),
   821 => (x"c7",x"c4",x"31",x"c4"),
   822 => (x"4b",x"26",x"59",x"f0"),
   823 => (x"c4",x"1e",x"4f",x"26"),
   824 => (x"49",x"bf",x"cc",x"cc"),
   825 => (x"bf",x"c0",x"cc",x"c4"),
   826 => (x"87",x"c4",x"05",x"a9"),
   827 => (x"87",x"c2",x"4a",x"c0"),
   828 => (x"48",x"72",x"4a",x"71"),
   829 => (x"5e",x"0e",x"4f",x"26"),
   830 => (x"71",x"0e",x"5c",x"5b"),
   831 => (x"72",x"4b",x"c0",x"4a"),
   832 => (x"e1",x"c0",x"02",x"9a"),
   833 => (x"49",x"a2",x"da",x"87"),
   834 => (x"c4",x"4b",x"69",x"9f"),
   835 => (x"02",x"bf",x"e8",x"c7"),
   836 => (x"a2",x"d4",x"87",x"cf"),
   837 => (x"49",x"69",x"9f",x"49"),
   838 => (x"ff",x"ff",x"c0",x"4c"),
   839 => (x"c2",x"34",x"d0",x"9c"),
   840 => (x"74",x"4c",x"c0",x"87"),
   841 => (x"49",x"73",x"b3",x"49"),
   842 => (x"26",x"87",x"d4",x"fd"),
   843 => (x"26",x"4b",x"26",x"4c"),
   844 => (x"5b",x"5e",x"0e",x"4f"),
   845 => (x"f0",x"0e",x"5d",x"5c"),
   846 => (x"59",x"a6",x"c8",x"86"),
   847 => (x"ff",x"ff",x"ff",x"cf"),
   848 => (x"7e",x"c0",x"4c",x"f8"),
   849 => (x"d8",x"02",x"66",x"c4"),
   850 => (x"dc",x"ff",x"c3",x"87"),
   851 => (x"c3",x"78",x"c0",x"48"),
   852 => (x"c4",x"48",x"d4",x"ff"),
   853 => (x"78",x"bf",x"d0",x"cc"),
   854 => (x"48",x"d8",x"ff",x"c3"),
   855 => (x"bf",x"cc",x"cc",x"c4"),
   856 => (x"fd",x"c7",x"c4",x"78"),
   857 => (x"c4",x"50",x"c0",x"48"),
   858 => (x"49",x"bf",x"ec",x"c7"),
   859 => (x"bf",x"dc",x"ff",x"c3"),
   860 => (x"03",x"aa",x"71",x"4a"),
   861 => (x"72",x"87",x"cc",x"c4"),
   862 => (x"05",x"99",x"cf",x"49"),
   863 => (x"c1",x"87",x"ea",x"c0"),
   864 => (x"c3",x"48",x"cc",x"c2"),
   865 => (x"78",x"bf",x"d4",x"ff"),
   866 => (x"1e",x"e0",x"ff",x"c3"),
   867 => (x"bf",x"d4",x"ff",x"c3"),
   868 => (x"d4",x"ff",x"c3",x"49"),
   869 => (x"78",x"a1",x"c1",x"48"),
   870 => (x"e1",x"dc",x"ff",x"71"),
   871 => (x"c0",x"86",x"c4",x"87"),
   872 => (x"c3",x"48",x"e8",x"fc"),
   873 => (x"cc",x"78",x"e0",x"ff"),
   874 => (x"e8",x"fc",x"c0",x"87"),
   875 => (x"e0",x"c0",x"48",x"bf"),
   876 => (x"ec",x"fc",x"c0",x"80"),
   877 => (x"dc",x"ff",x"c3",x"58"),
   878 => (x"80",x"c1",x"48",x"bf"),
   879 => (x"58",x"e0",x"ff",x"c3"),
   880 => (x"00",x"0f",x"28",x"27"),
   881 => (x"bf",x"97",x"bf",x"00"),
   882 => (x"c2",x"02",x"9d",x"4d"),
   883 => (x"e5",x"c3",x"87",x"e5"),
   884 => (x"de",x"c2",x"02",x"ad"),
   885 => (x"e8",x"fc",x"c0",x"87"),
   886 => (x"a3",x"cb",x"4b",x"bf"),
   887 => (x"cf",x"4c",x"11",x"49"),
   888 => (x"d2",x"c1",x"05",x"ac"),
   889 => (x"df",x"49",x"75",x"87"),
   890 => (x"cd",x"89",x"c1",x"99"),
   891 => (x"f0",x"c7",x"c4",x"91"),
   892 => (x"4a",x"a3",x"c1",x"81"),
   893 => (x"a3",x"c3",x"51",x"12"),
   894 => (x"c5",x"51",x"12",x"4a"),
   895 => (x"51",x"12",x"4a",x"a3"),
   896 => (x"12",x"4a",x"a3",x"c7"),
   897 => (x"4a",x"a3",x"c9",x"51"),
   898 => (x"a3",x"ce",x"51",x"12"),
   899 => (x"d0",x"51",x"12",x"4a"),
   900 => (x"51",x"12",x"4a",x"a3"),
   901 => (x"12",x"4a",x"a3",x"d2"),
   902 => (x"4a",x"a3",x"d4",x"51"),
   903 => (x"a3",x"d6",x"51",x"12"),
   904 => (x"d8",x"51",x"12",x"4a"),
   905 => (x"51",x"12",x"4a",x"a3"),
   906 => (x"12",x"4a",x"a3",x"dc"),
   907 => (x"4a",x"a3",x"de",x"51"),
   908 => (x"7e",x"c1",x"51",x"12"),
   909 => (x"74",x"87",x"fc",x"c0"),
   910 => (x"05",x"99",x"c8",x"49"),
   911 => (x"74",x"87",x"ed",x"c0"),
   912 => (x"05",x"99",x"d0",x"49"),
   913 => (x"e0",x"c0",x"87",x"d3"),
   914 => (x"cc",x"c0",x"02",x"66"),
   915 => (x"c0",x"49",x"73",x"87"),
   916 => (x"70",x"0f",x"66",x"e0"),
   917 => (x"d3",x"c0",x"02",x"98"),
   918 => (x"c0",x"05",x"6e",x"87"),
   919 => (x"c7",x"c4",x"87",x"c6"),
   920 => (x"50",x"c0",x"48",x"f0"),
   921 => (x"bf",x"e8",x"fc",x"c0"),
   922 => (x"87",x"eb",x"c2",x"48"),
   923 => (x"48",x"fd",x"c7",x"c4"),
   924 => (x"c4",x"7e",x"50",x"c0"),
   925 => (x"49",x"bf",x"ec",x"c7"),
   926 => (x"bf",x"dc",x"ff",x"c3"),
   927 => (x"04",x"aa",x"71",x"4a"),
   928 => (x"cf",x"87",x"f4",x"fb"),
   929 => (x"f8",x"ff",x"ff",x"ff"),
   930 => (x"d0",x"cc",x"c4",x"4c"),
   931 => (x"c8",x"c0",x"05",x"bf"),
   932 => (x"e8",x"c7",x"c4",x"87"),
   933 => (x"fc",x"c1",x"02",x"bf"),
   934 => (x"d8",x"ff",x"c3",x"87"),
   935 => (x"db",x"e6",x"49",x"bf"),
   936 => (x"dc",x"ff",x"c3",x"87"),
   937 => (x"48",x"a6",x"c4",x"58"),
   938 => (x"bf",x"d8",x"ff",x"c3"),
   939 => (x"e8",x"c7",x"c4",x"78"),
   940 => (x"db",x"c0",x"02",x"bf"),
   941 => (x"49",x"66",x"c4",x"87"),
   942 => (x"a9",x"74",x"99",x"74"),
   943 => (x"87",x"c8",x"c0",x"02"),
   944 => (x"c0",x"48",x"a6",x"c8"),
   945 => (x"87",x"e7",x"c0",x"78"),
   946 => (x"c1",x"48",x"a6",x"c8"),
   947 => (x"87",x"df",x"c0",x"78"),
   948 => (x"cf",x"49",x"66",x"c4"),
   949 => (x"a9",x"99",x"f8",x"ff"),
   950 => (x"87",x"c8",x"c0",x"02"),
   951 => (x"c0",x"48",x"a6",x"cc"),
   952 => (x"87",x"c5",x"c0",x"78"),
   953 => (x"c1",x"48",x"a6",x"cc"),
   954 => (x"48",x"a6",x"c8",x"78"),
   955 => (x"c8",x"78",x"66",x"cc"),
   956 => (x"e0",x"c0",x"05",x"66"),
   957 => (x"49",x"66",x"c4",x"87"),
   958 => (x"c7",x"c4",x"89",x"c2"),
   959 => (x"91",x"4a",x"bf",x"e0"),
   960 => (x"bf",x"fc",x"cb",x"c4"),
   961 => (x"d4",x"ff",x"c3",x"4a"),
   962 => (x"78",x"a1",x"72",x"48"),
   963 => (x"48",x"dc",x"ff",x"c3"),
   964 => (x"d2",x"f9",x"78",x"c0"),
   965 => (x"cf",x"48",x"c0",x"87"),
   966 => (x"f8",x"ff",x"ff",x"ff"),
   967 => (x"26",x"8e",x"f0",x"4c"),
   968 => (x"26",x"4c",x"26",x"4d"),
   969 => (x"00",x"4f",x"26",x"4b"),
   970 => (x"00",x"00",x"00",x"00"),
   971 => (x"5c",x"5b",x"5e",x"0e"),
   972 => (x"86",x"fc",x"0e",x"5d"),
   973 => (x"49",x"6e",x"7e",x"71"),
   974 => (x"c0",x"87",x"c4",x"f5"),
   975 => (x"49",x"49",x"c1",x"1e"),
   976 => (x"c4",x"87",x"ee",x"f7"),
   977 => (x"9a",x"4a",x"70",x"86"),
   978 => (x"87",x"c7",x"c1",x"02"),
   979 => (x"9f",x"49",x"a2",x"da"),
   980 => (x"c7",x"c4",x"4b",x"69"),
   981 => (x"cf",x"02",x"bf",x"e8"),
   982 => (x"49",x"a2",x"d4",x"87"),
   983 => (x"4c",x"49",x"69",x"9f"),
   984 => (x"9c",x"ff",x"ff",x"c0"),
   985 => (x"87",x"c2",x"34",x"d0"),
   986 => (x"49",x"74",x"4c",x"c0"),
   987 => (x"66",x"d4",x"4b",x"a3"),
   988 => (x"87",x"c4",x"05",x"ab"),
   989 => (x"87",x"dd",x"48",x"c1"),
   990 => (x"9a",x"72",x"1e",x"c0"),
   991 => (x"c0",x"87",x"c4",x"02"),
   992 => (x"c1",x"87",x"c2",x"4d"),
   993 => (x"f6",x"49",x"75",x"4d"),
   994 => (x"86",x"c4",x"87",x"e7"),
   995 => (x"05",x"9a",x"4a",x"70"),
   996 => (x"c0",x"87",x"f9",x"fe"),
   997 => (x"26",x"8e",x"fc",x"48"),
   998 => (x"26",x"4c",x"26",x"4d"),
   999 => (x"0e",x"4f",x"26",x"4b"),
  1000 => (x"5d",x"5c",x"5b",x"5e"),
  1001 => (x"c8",x"86",x"f4",x"0e"),
  1002 => (x"66",x"c4",x"59",x"a6"),
  1003 => (x"48",x"87",x"c9",x"02"),
  1004 => (x"bf",x"c0",x"cc",x"c4"),
  1005 => (x"87",x"c5",x"05",x"a8"),
  1006 => (x"f9",x"c2",x"48",x"c1"),
  1007 => (x"49",x"66",x"c4",x"87"),
  1008 => (x"c7",x"c4",x"89",x"c2"),
  1009 => (x"91",x"4a",x"bf",x"e0"),
  1010 => (x"bf",x"fc",x"cb",x"c4"),
  1011 => (x"c3",x"49",x"a1",x"4a"),
  1012 => (x"71",x"1e",x"e0",x"ff"),
  1013 => (x"87",x"e6",x"d3",x"ff"),
  1014 => (x"98",x"70",x"86",x"c4"),
  1015 => (x"c0",x"87",x"c5",x"05"),
  1016 => (x"87",x"d2",x"c2",x"48"),
  1017 => (x"4c",x"e0",x"ff",x"c3"),
  1018 => (x"6c",x"97",x"7e",x"c0"),
  1019 => (x"58",x"a6",x"cc",x"48"),
  1020 => (x"c1",x"02",x"98",x"70"),
  1021 => (x"c3",x"48",x"87",x"ee"),
  1022 => (x"c1",x"02",x"a8",x"e5"),
  1023 => (x"a4",x"cb",x"87",x"e6"),
  1024 => (x"49",x"69",x"97",x"49"),
  1025 => (x"c1",x"02",x"99",x"d0"),
  1026 => (x"4a",x"74",x"87",x"da"),
  1027 => (x"49",x"c0",x"c2",x"c1"),
  1028 => (x"c1",x"ff",x"4b",x"c8"),
  1029 => (x"98",x"70",x"87",x"ee"),
  1030 => (x"87",x"c8",x"c1",x"05"),
  1031 => (x"c4",x"7e",x"a4",x"da"),
  1032 => (x"02",x"bf",x"e8",x"c7"),
  1033 => (x"a4",x"d4",x"87",x"cf"),
  1034 => (x"49",x"69",x"9f",x"49"),
  1035 => (x"ff",x"ff",x"c0",x"4d"),
  1036 => (x"c2",x"35",x"d0",x"9d"),
  1037 => (x"6e",x"4d",x"c0",x"87"),
  1038 => (x"c8",x"49",x"bf",x"9f"),
  1039 => (x"a5",x"71",x"48",x"a6"),
  1040 => (x"da",x"fd",x"49",x"78"),
  1041 => (x"02",x"98",x"70",x"87"),
  1042 => (x"66",x"c4",x"87",x"d4"),
  1043 => (x"49",x"66",x"cc",x"1e"),
  1044 => (x"c4",x"87",x"d9",x"fb"),
  1045 => (x"02",x"98",x"70",x"86"),
  1046 => (x"7e",x"c1",x"87",x"c4"),
  1047 => (x"7e",x"c0",x"87",x"c2"),
  1048 => (x"87",x"d2",x"48",x"6e"),
  1049 => (x"6e",x"84",x"e0",x"c0"),
  1050 => (x"70",x"80",x"c1",x"48"),
  1051 => (x"a8",x"d0",x"48",x"7e"),
  1052 => (x"87",x"f6",x"fd",x"04"),
  1053 => (x"8e",x"f4",x"48",x"c0"),
  1054 => (x"4c",x"26",x"4d",x"26"),
  1055 => (x"4f",x"26",x"4b",x"26"),
  1056 => (x"20",x"20",x"2e",x"2e"),
  1057 => (x"20",x"20",x"20",x"20"),
  1058 => (x"00",x"20",x"20",x"20"),
  1059 => (x"ff",x"ff",x"ff",x"ff"),
  1060 => (x"00",x"00",x"10",x"98"),
  1061 => (x"00",x"00",x"10",x"a4"),
  1062 => (x"33",x"54",x"41",x"46"),
  1063 => (x"20",x"20",x"20",x"32"),
  1064 => (x"00",x"00",x"00",x"00"),
  1065 => (x"31",x"54",x"41",x"46"),
  1066 => (x"20",x"20",x"20",x"36"),
  1067 => (x"d0",x"ff",x"1e",x"00"),
  1068 => (x"78",x"e0",x"c0",x"48"),
  1069 => (x"c2",x"1e",x"4f",x"26"),
  1070 => (x"70",x"87",x"dd",x"d2"),
  1071 => (x"c6",x"02",x"99",x"49"),
  1072 => (x"a9",x"fb",x"c0",x"87"),
  1073 => (x"71",x"87",x"f0",x"05"),
  1074 => (x"0e",x"4f",x"26",x"48"),
  1075 => (x"0e",x"5c",x"5b",x"5e"),
  1076 => (x"4c",x"c0",x"4b",x"71"),
  1077 => (x"87",x"c0",x"d2",x"c2"),
  1078 => (x"02",x"99",x"49",x"70"),
  1079 => (x"c0",x"87",x"fa",x"c0"),
  1080 => (x"c0",x"02",x"a9",x"ec"),
  1081 => (x"fb",x"c0",x"87",x"f3"),
  1082 => (x"ec",x"c0",x"02",x"a9"),
  1083 => (x"b7",x"66",x"cc",x"87"),
  1084 => (x"87",x"c7",x"03",x"ac"),
  1085 => (x"c2",x"02",x"66",x"d0"),
  1086 => (x"71",x"53",x"71",x"87"),
  1087 => (x"87",x"c2",x"02",x"99"),
  1088 => (x"d1",x"c2",x"84",x"c1"),
  1089 => (x"49",x"70",x"87",x"d2"),
  1090 => (x"87",x"cd",x"02",x"99"),
  1091 => (x"02",x"a9",x"ec",x"c0"),
  1092 => (x"fb",x"c0",x"87",x"c7"),
  1093 => (x"d4",x"ff",x"05",x"a9"),
  1094 => (x"02",x"66",x"d0",x"87"),
  1095 => (x"97",x"c0",x"87",x"c3"),
  1096 => (x"a9",x"ec",x"c0",x"7b"),
  1097 => (x"74",x"87",x"c4",x"05"),
  1098 => (x"74",x"87",x"c5",x"4a"),
  1099 => (x"8a",x"0a",x"c0",x"4a"),
  1100 => (x"4c",x"26",x"48",x"72"),
  1101 => (x"4f",x"26",x"4b",x"26"),
  1102 => (x"db",x"d0",x"c2",x"1e"),
  1103 => (x"c0",x"4a",x"70",x"87"),
  1104 => (x"c9",x"04",x"aa",x"f0"),
  1105 => (x"aa",x"f9",x"c0",x"87"),
  1106 => (x"c0",x"87",x"c3",x"01"),
  1107 => (x"c1",x"c1",x"8a",x"f0"),
  1108 => (x"87",x"c9",x"04",x"aa"),
  1109 => (x"01",x"aa",x"da",x"c1"),
  1110 => (x"f7",x"c0",x"87",x"c3"),
  1111 => (x"26",x"48",x"72",x"8a"),
  1112 => (x"5b",x"5e",x"0e",x"4f"),
  1113 => (x"f8",x"0e",x"5d",x"5c"),
  1114 => (x"c0",x"4c",x"71",x"86"),
  1115 => (x"ca",x"d0",x"c2",x"7e"),
  1116 => (x"c1",x"4b",x"c0",x"87"),
  1117 => (x"bf",x"97",x"c4",x"c8"),
  1118 => (x"04",x"a9",x"c0",x"49"),
  1119 => (x"f5",x"fc",x"87",x"cf"),
  1120 => (x"c1",x"83",x"c1",x"87"),
  1121 => (x"bf",x"97",x"c4",x"c8"),
  1122 => (x"f1",x"06",x"ab",x"49"),
  1123 => (x"c4",x"c8",x"c1",x"87"),
  1124 => (x"d0",x"02",x"bf",x"97"),
  1125 => (x"ff",x"ce",x"c2",x"87"),
  1126 => (x"99",x"49",x"70",x"87"),
  1127 => (x"c0",x"87",x"c6",x"02"),
  1128 => (x"f0",x"05",x"a9",x"ec"),
  1129 => (x"c2",x"4b",x"c0",x"87"),
  1130 => (x"70",x"87",x"ed",x"ce"),
  1131 => (x"e7",x"ce",x"c2",x"4d"),
  1132 => (x"58",x"a6",x"c8",x"87"),
  1133 => (x"87",x"e0",x"ce",x"c2"),
  1134 => (x"83",x"c1",x"4a",x"70"),
  1135 => (x"97",x"49",x"a4",x"c8"),
  1136 => (x"05",x"ad",x"49",x"69"),
  1137 => (x"a4",x"c9",x"87",x"da"),
  1138 => (x"49",x"69",x"97",x"49"),
  1139 => (x"05",x"a9",x"66",x"c4"),
  1140 => (x"a4",x"ca",x"87",x"ce"),
  1141 => (x"49",x"69",x"97",x"49"),
  1142 => (x"87",x"c4",x"05",x"aa"),
  1143 => (x"87",x"d0",x"7e",x"c1"),
  1144 => (x"02",x"ad",x"ec",x"c0"),
  1145 => (x"fb",x"c0",x"87",x"c6"),
  1146 => (x"87",x"c4",x"05",x"ad"),
  1147 => (x"7e",x"c1",x"4b",x"c0"),
  1148 => (x"f2",x"fe",x"02",x"6e"),
  1149 => (x"87",x"f5",x"fa",x"87"),
  1150 => (x"8e",x"f8",x"48",x"73"),
  1151 => (x"4c",x"26",x"4d",x"26"),
  1152 => (x"4f",x"26",x"4b",x"26"),
  1153 => (x"5b",x"5e",x"0e",x"00"),
  1154 => (x"f4",x"0e",x"5d",x"5c"),
  1155 => (x"ff",x"7e",x"71",x"86"),
  1156 => (x"1e",x"6e",x"4b",x"d4"),
  1157 => (x"49",x"dc",x"cc",x"c4"),
  1158 => (x"87",x"d7",x"da",x"ff"),
  1159 => (x"98",x"70",x"86",x"c4"),
  1160 => (x"87",x"f7",x"c4",x"02"),
  1161 => (x"c1",x"48",x"a6",x"c4"),
  1162 => (x"78",x"bf",x"e8",x"f3"),
  1163 => (x"f0",x"fc",x"49",x"6e"),
  1164 => (x"58",x"a6",x"cc",x"87"),
  1165 => (x"c5",x"05",x"98",x"70"),
  1166 => (x"48",x"a6",x"c8",x"87"),
  1167 => (x"d0",x"ff",x"78",x"c1"),
  1168 => (x"c1",x"78",x"c5",x"48"),
  1169 => (x"66",x"c8",x"7b",x"d5"),
  1170 => (x"c6",x"89",x"c1",x"49"),
  1171 => (x"e0",x"f3",x"c1",x"31"),
  1172 => (x"48",x"4a",x"bf",x"97"),
  1173 => (x"7b",x"70",x"b0",x"71"),
  1174 => (x"c4",x"48",x"d0",x"ff"),
  1175 => (x"d4",x"cc",x"c4",x"78"),
  1176 => (x"d0",x"49",x"bf",x"97"),
  1177 => (x"87",x"d7",x"02",x"99"),
  1178 => (x"d6",x"c1",x"78",x"c5"),
  1179 => (x"c3",x"4a",x"c0",x"7b"),
  1180 => (x"82",x"c1",x"7b",x"ff"),
  1181 => (x"04",x"aa",x"e0",x"c0"),
  1182 => (x"d0",x"ff",x"87",x"f5"),
  1183 => (x"c3",x"78",x"c4",x"48"),
  1184 => (x"d0",x"ff",x"7b",x"ff"),
  1185 => (x"c1",x"78",x"c5",x"48"),
  1186 => (x"7b",x"c1",x"7b",x"d3"),
  1187 => (x"7e",x"73",x"78",x"c4"),
  1188 => (x"c0",x"48",x"66",x"c4"),
  1189 => (x"c2",x"06",x"a8",x"b7"),
  1190 => (x"cc",x"c4",x"87",x"ee"),
  1191 => (x"c4",x"4c",x"bf",x"e4"),
  1192 => (x"88",x"74",x"48",x"66"),
  1193 => (x"74",x"58",x"a6",x"c8"),
  1194 => (x"f7",x"c1",x"02",x"9c"),
  1195 => (x"e0",x"ff",x"c3",x"87"),
  1196 => (x"4b",x"c0",x"c8",x"4d"),
  1197 => (x"ac",x"b7",x"c0",x"8c"),
  1198 => (x"c8",x"87",x"c6",x"03"),
  1199 => (x"c0",x"4b",x"a4",x"c0"),
  1200 => (x"d4",x"cc",x"c4",x"4c"),
  1201 => (x"d0",x"49",x"bf",x"97"),
  1202 => (x"87",x"d1",x"02",x"99"),
  1203 => (x"cc",x"c4",x"1e",x"c0"),
  1204 => (x"dd",x"ff",x"49",x"dc"),
  1205 => (x"86",x"c4",x"87",x"e1"),
  1206 => (x"eb",x"c0",x"4a",x"70"),
  1207 => (x"e0",x"ff",x"c3",x"87"),
  1208 => (x"dc",x"cc",x"c4",x"1e"),
  1209 => (x"ce",x"dd",x"ff",x"49"),
  1210 => (x"70",x"86",x"c4",x"87"),
  1211 => (x"48",x"d0",x"ff",x"4a"),
  1212 => (x"6e",x"78",x"c5",x"c8"),
  1213 => (x"78",x"d4",x"c1",x"48"),
  1214 => (x"08",x"6e",x"48",x"15"),
  1215 => (x"05",x"8b",x"c1",x"78"),
  1216 => (x"ff",x"87",x"f5",x"ff"),
  1217 => (x"78",x"c4",x"48",x"d0"),
  1218 => (x"c5",x"05",x"9a",x"72"),
  1219 => (x"c1",x"48",x"c0",x"87"),
  1220 => (x"1e",x"c1",x"87",x"cb"),
  1221 => (x"49",x"dc",x"cc",x"c4"),
  1222 => (x"87",x"fb",x"da",x"ff"),
  1223 => (x"9c",x"74",x"86",x"c4"),
  1224 => (x"87",x"c9",x"fe",x"05"),
  1225 => (x"c0",x"48",x"66",x"c4"),
  1226 => (x"d1",x"06",x"a8",x"b7"),
  1227 => (x"dc",x"cc",x"c4",x"87"),
  1228 => (x"d0",x"78",x"c0",x"48"),
  1229 => (x"f4",x"78",x"c0",x"80"),
  1230 => (x"e8",x"cc",x"c4",x"80"),
  1231 => (x"66",x"c4",x"78",x"bf"),
  1232 => (x"a8",x"b7",x"c0",x"48"),
  1233 => (x"87",x"d2",x"fd",x"01"),
  1234 => (x"d0",x"ff",x"4b",x"6e"),
  1235 => (x"c1",x"78",x"c5",x"48"),
  1236 => (x"7b",x"c0",x"7b",x"d3"),
  1237 => (x"48",x"c1",x"78",x"c4"),
  1238 => (x"c0",x"87",x"c2",x"c0"),
  1239 => (x"26",x"8e",x"f4",x"48"),
  1240 => (x"26",x"4c",x"26",x"4d"),
  1241 => (x"0e",x"4f",x"26",x"4b"),
  1242 => (x"5d",x"5c",x"5b",x"5e"),
  1243 => (x"71",x"86",x"fc",x"0e"),
  1244 => (x"4c",x"4b",x"c0",x"4d"),
  1245 => (x"e8",x"c0",x"04",x"ad"),
  1246 => (x"e1",x"c5",x"c1",x"87"),
  1247 => (x"02",x"9c",x"74",x"1e"),
  1248 => (x"4a",x"c0",x"87",x"c4"),
  1249 => (x"4a",x"c1",x"87",x"c2"),
  1250 => (x"e4",x"e6",x"49",x"72"),
  1251 => (x"70",x"86",x"c4",x"87"),
  1252 => (x"6e",x"83",x"c1",x"7e"),
  1253 => (x"75",x"87",x"c2",x"05"),
  1254 => (x"75",x"84",x"c1",x"4b"),
  1255 => (x"d8",x"ff",x"06",x"ab"),
  1256 => (x"fc",x"48",x"6e",x"87"),
  1257 => (x"26",x"4d",x"26",x"8e"),
  1258 => (x"26",x"4b",x"26",x"4c"),
  1259 => (x"5b",x"5e",x"0e",x"4f"),
  1260 => (x"fc",x"0e",x"5d",x"5c"),
  1261 => (x"49",x"4c",x"71",x"86"),
  1262 => (x"cd",x"c4",x"91",x"de"),
  1263 => (x"85",x"71",x"4d",x"f8"),
  1264 => (x"c1",x"02",x"6d",x"97"),
  1265 => (x"cd",x"c4",x"87",x"dd"),
  1266 => (x"74",x"49",x"bf",x"e4"),
  1267 => (x"d6",x"fe",x"71",x"81"),
  1268 => (x"48",x"7e",x"70",x"87"),
  1269 => (x"f3",x"c0",x"02",x"98"),
  1270 => (x"ec",x"cd",x"c4",x"87"),
  1271 => (x"cb",x"4a",x"70",x"4b"),
  1272 => (x"dd",x"f3",x"fe",x"49"),
  1273 => (x"cc",x"4b",x"74",x"87"),
  1274 => (x"fc",x"f3",x"c1",x"93"),
  1275 => (x"c1",x"83",x"c4",x"83"),
  1276 => (x"74",x"7b",x"f0",x"d0"),
  1277 => (x"e7",x"c6",x"c1",x"49"),
  1278 => (x"c1",x"7b",x"75",x"87"),
  1279 => (x"bf",x"97",x"e4",x"f3"),
  1280 => (x"cd",x"c4",x"1e",x"49"),
  1281 => (x"d5",x"c2",x"49",x"ec"),
  1282 => (x"86",x"c4",x"87",x"d6"),
  1283 => (x"c6",x"c1",x"49",x"74"),
  1284 => (x"49",x"c0",x"87",x"ce"),
  1285 => (x"87",x"e9",x"c7",x"c1"),
  1286 => (x"48",x"d8",x"cc",x"c4"),
  1287 => (x"49",x"c1",x"78",x"c0"),
  1288 => (x"fc",x"87",x"c4",x"de"),
  1289 => (x"26",x"4d",x"26",x"8e"),
  1290 => (x"26",x"4b",x"26",x"4c"),
  1291 => (x"00",x"00",x"00",x"4f"),
  1292 => (x"64",x"61",x"6f",x"4c"),
  1293 => (x"2e",x"67",x"6e",x"69"),
  1294 => (x"1e",x"00",x"2e",x"2e"),
  1295 => (x"4a",x"71",x"1e",x"73"),
  1296 => (x"e4",x"cd",x"c4",x"49"),
  1297 => (x"fc",x"71",x"81",x"bf"),
  1298 => (x"4b",x"70",x"87",x"dd"),
  1299 => (x"87",x"c4",x"02",x"9b"),
  1300 => (x"87",x"e2",x"e2",x"49"),
  1301 => (x"48",x"e4",x"cd",x"c4"),
  1302 => (x"49",x"c1",x"78",x"c0"),
  1303 => (x"26",x"87",x"c8",x"dd"),
  1304 => (x"1e",x"4f",x"26",x"4b"),
  1305 => (x"c6",x"c1",x"49",x"c0"),
  1306 => (x"4f",x"26",x"87",x"d7"),
  1307 => (x"49",x"4a",x"71",x"1e"),
  1308 => (x"f3",x"c1",x"91",x"cc"),
  1309 => (x"81",x"c8",x"81",x"fc"),
  1310 => (x"cc",x"c4",x"48",x"11"),
  1311 => (x"cd",x"c4",x"58",x"dc"),
  1312 => (x"78",x"c0",x"48",x"e4"),
  1313 => (x"de",x"dc",x"49",x"c1"),
  1314 => (x"1e",x"4f",x"26",x"87"),
  1315 => (x"d2",x"02",x"99",x"71"),
  1316 => (x"d8",x"f5",x"c1",x"87"),
  1317 => (x"f7",x"50",x"c0",x"48"),
  1318 => (x"ec",x"d1",x"c1",x"80"),
  1319 => (x"f4",x"f3",x"c1",x"40"),
  1320 => (x"c1",x"87",x"ce",x"78"),
  1321 => (x"c1",x"48",x"d4",x"f5"),
  1322 => (x"fc",x"78",x"ec",x"f3"),
  1323 => (x"e3",x"d1",x"c1",x"80"),
  1324 => (x"0e",x"4f",x"26",x"78"),
  1325 => (x"5d",x"5c",x"5b",x"5e"),
  1326 => (x"c3",x"86",x"f4",x"0e"),
  1327 => (x"c0",x"4d",x"e0",x"ff"),
  1328 => (x"48",x"a6",x"c8",x"4c"),
  1329 => (x"7e",x"75",x"78",x"c0"),
  1330 => (x"bf",x"e4",x"cd",x"c4"),
  1331 => (x"06",x"a8",x"c0",x"48"),
  1332 => (x"c8",x"87",x"c0",x"c1"),
  1333 => (x"7e",x"75",x"5c",x"a6"),
  1334 => (x"48",x"e0",x"ff",x"c3"),
  1335 => (x"f2",x"c0",x"02",x"98"),
  1336 => (x"4d",x"66",x"c4",x"87"),
  1337 => (x"1e",x"e1",x"c5",x"c1"),
  1338 => (x"c4",x"02",x"66",x"cc"),
  1339 => (x"c2",x"4c",x"c0",x"87"),
  1340 => (x"74",x"4c",x"c1",x"87"),
  1341 => (x"87",x"f9",x"e0",x"49"),
  1342 => (x"7e",x"70",x"86",x"c4"),
  1343 => (x"66",x"c8",x"85",x"c1"),
  1344 => (x"cc",x"80",x"c1",x"48"),
  1345 => (x"cd",x"c4",x"58",x"a6"),
  1346 => (x"03",x"ad",x"bf",x"e4"),
  1347 => (x"05",x"6e",x"87",x"c5"),
  1348 => (x"6e",x"87",x"d1",x"ff"),
  1349 => (x"75",x"4c",x"c0",x"4d"),
  1350 => (x"dd",x"c3",x"02",x"9d"),
  1351 => (x"e1",x"c5",x"c1",x"87"),
  1352 => (x"02",x"66",x"cc",x"1e"),
  1353 => (x"a6",x"c8",x"87",x"c7"),
  1354 => (x"c5",x"78",x"c0",x"48"),
  1355 => (x"48",x"a6",x"c8",x"87"),
  1356 => (x"66",x"c8",x"78",x"c1"),
  1357 => (x"f8",x"df",x"ff",x"49"),
  1358 => (x"70",x"86",x"c4",x"87"),
  1359 => (x"02",x"98",x"48",x"7e"),
  1360 => (x"49",x"87",x"e4",x"c2"),
  1361 => (x"69",x"97",x"81",x"cb"),
  1362 => (x"02",x"99",x"d0",x"49"),
  1363 => (x"74",x"87",x"d4",x"c1"),
  1364 => (x"c1",x"91",x"cc",x"49"),
  1365 => (x"c1",x"81",x"fc",x"f3"),
  1366 => (x"c8",x"79",x"fb",x"d0"),
  1367 => (x"51",x"ff",x"c3",x"81"),
  1368 => (x"91",x"de",x"49",x"74"),
  1369 => (x"4d",x"f8",x"cd",x"c4"),
  1370 => (x"c1",x"c2",x"85",x"71"),
  1371 => (x"a5",x"c1",x"7d",x"97"),
  1372 => (x"51",x"e0",x"c0",x"49"),
  1373 => (x"97",x"f0",x"c7",x"c4"),
  1374 => (x"87",x"d2",x"02",x"bf"),
  1375 => (x"a5",x"c2",x"84",x"c1"),
  1376 => (x"f0",x"c7",x"c4",x"4b"),
  1377 => (x"fe",x"49",x"db",x"4a"),
  1378 => (x"c1",x"87",x"f7",x"ec"),
  1379 => (x"a5",x"cd",x"87",x"d9"),
  1380 => (x"c1",x"51",x"c0",x"49"),
  1381 => (x"4b",x"a5",x"c2",x"84"),
  1382 => (x"49",x"cb",x"4a",x"6e"),
  1383 => (x"87",x"e2",x"ec",x"fe"),
  1384 => (x"74",x"87",x"c4",x"c1"),
  1385 => (x"c1",x"91",x"cc",x"49"),
  1386 => (x"c1",x"81",x"fc",x"f3"),
  1387 => (x"c4",x"79",x"ed",x"ce"),
  1388 => (x"bf",x"97",x"f0",x"c7"),
  1389 => (x"74",x"87",x"d8",x"02"),
  1390 => (x"c1",x"91",x"de",x"49"),
  1391 => (x"f8",x"cd",x"c4",x"84"),
  1392 => (x"c4",x"83",x"71",x"4b"),
  1393 => (x"dd",x"4a",x"f0",x"c7"),
  1394 => (x"f5",x"eb",x"fe",x"49"),
  1395 => (x"74",x"87",x"d8",x"87"),
  1396 => (x"c4",x"93",x"de",x"4b"),
  1397 => (x"cb",x"83",x"f8",x"cd"),
  1398 => (x"51",x"c0",x"49",x"a3"),
  1399 => (x"6e",x"73",x"84",x"c1"),
  1400 => (x"fe",x"49",x"cb",x"4a"),
  1401 => (x"c8",x"87",x"db",x"eb"),
  1402 => (x"80",x"c1",x"48",x"66"),
  1403 => (x"c7",x"58",x"a6",x"cc"),
  1404 => (x"c5",x"c0",x"03",x"ac"),
  1405 => (x"fc",x"05",x"6e",x"87"),
  1406 => (x"48",x"74",x"87",x"e3"),
  1407 => (x"4d",x"26",x"8e",x"f4"),
  1408 => (x"4b",x"26",x"4c",x"26"),
  1409 => (x"73",x"1e",x"4f",x"26"),
  1410 => (x"49",x"4b",x"71",x"1e"),
  1411 => (x"f3",x"c1",x"91",x"cc"),
  1412 => (x"a1",x"c8",x"81",x"fc"),
  1413 => (x"e0",x"f3",x"c1",x"4a"),
  1414 => (x"c9",x"50",x"12",x"48"),
  1415 => (x"c8",x"c1",x"4a",x"a1"),
  1416 => (x"50",x"12",x"48",x"c4"),
  1417 => (x"f3",x"c1",x"81",x"ca"),
  1418 => (x"50",x"11",x"48",x"e4"),
  1419 => (x"97",x"e4",x"f3",x"c1"),
  1420 => (x"c0",x"1e",x"49",x"bf"),
  1421 => (x"e7",x"cc",x"c2",x"49"),
  1422 => (x"d8",x"cc",x"c4",x"87"),
  1423 => (x"c1",x"78",x"de",x"48"),
  1424 => (x"87",x"e3",x"d5",x"49"),
  1425 => (x"4b",x"26",x"8e",x"fc"),
  1426 => (x"5e",x"0e",x"4f",x"26"),
  1427 => (x"0e",x"5d",x"5c",x"5b"),
  1428 => (x"4d",x"71",x"86",x"f4"),
  1429 => (x"c1",x"91",x"cc",x"49"),
  1430 => (x"c8",x"81",x"fc",x"f3"),
  1431 => (x"a1",x"ca",x"4a",x"a1"),
  1432 => (x"48",x"a6",x"c4",x"7e"),
  1433 => (x"bf",x"f4",x"d1",x"c4"),
  1434 => (x"bf",x"97",x"6e",x"78"),
  1435 => (x"4c",x"66",x"c4",x"4b"),
  1436 => (x"48",x"12",x"2c",x"73"),
  1437 => (x"70",x"58",x"a6",x"cc"),
  1438 => (x"c9",x"84",x"c1",x"9c"),
  1439 => (x"49",x"69",x"97",x"81"),
  1440 => (x"c2",x"04",x"ac",x"b7"),
  1441 => (x"6e",x"4c",x"c0",x"87"),
  1442 => (x"c8",x"4a",x"bf",x"97"),
  1443 => (x"31",x"72",x"49",x"66"),
  1444 => (x"66",x"c4",x"b9",x"ff"),
  1445 => (x"72",x"48",x"74",x"99"),
  1446 => (x"48",x"4a",x"70",x"30"),
  1447 => (x"d1",x"c4",x"b0",x"71"),
  1448 => (x"f9",x"c1",x"58",x"f8"),
  1449 => (x"49",x"c0",x"87",x"f9"),
  1450 => (x"75",x"87",x"fc",x"d3"),
  1451 => (x"ef",x"fb",x"c0",x"49"),
  1452 => (x"26",x"8e",x"f4",x"87"),
  1453 => (x"26",x"4c",x"26",x"4d"),
  1454 => (x"1e",x"4f",x"26",x"4b"),
  1455 => (x"4b",x"71",x"1e",x"73"),
  1456 => (x"02",x"4a",x"a3",x"c6"),
  1457 => (x"8a",x"c1",x"87",x"db"),
  1458 => (x"8a",x"87",x"d6",x"02"),
  1459 => (x"87",x"da",x"c1",x"02"),
  1460 => (x"fc",x"c0",x"02",x"8a"),
  1461 => (x"c0",x"02",x"8a",x"87"),
  1462 => (x"02",x"8a",x"87",x"e1"),
  1463 => (x"db",x"c1",x"87",x"cb"),
  1464 => (x"f6",x"49",x"c7",x"87"),
  1465 => (x"de",x"c1",x"87",x"c6"),
  1466 => (x"e4",x"cd",x"c4",x"87"),
  1467 => (x"cb",x"c1",x"02",x"bf"),
  1468 => (x"88",x"c1",x"48",x"87"),
  1469 => (x"58",x"e8",x"cd",x"c4"),
  1470 => (x"c4",x"87",x"c1",x"c1"),
  1471 => (x"02",x"bf",x"e8",x"cd"),
  1472 => (x"c4",x"87",x"f9",x"c0"),
  1473 => (x"48",x"bf",x"e4",x"cd"),
  1474 => (x"cd",x"c4",x"80",x"c1"),
  1475 => (x"eb",x"c0",x"58",x"e8"),
  1476 => (x"e4",x"cd",x"c4",x"87"),
  1477 => (x"89",x"c6",x"49",x"bf"),
  1478 => (x"59",x"e8",x"cd",x"c4"),
  1479 => (x"03",x"a9",x"b7",x"c0"),
  1480 => (x"cd",x"c4",x"87",x"da"),
  1481 => (x"78",x"c0",x"48",x"e4"),
  1482 => (x"cd",x"c4",x"87",x"d2"),
  1483 => (x"cb",x"02",x"bf",x"e8"),
  1484 => (x"e4",x"cd",x"c4",x"87"),
  1485 => (x"80",x"c6",x"48",x"bf"),
  1486 => (x"58",x"e8",x"cd",x"c4"),
  1487 => (x"e6",x"d1",x"49",x"c0"),
  1488 => (x"c0",x"49",x"73",x"87"),
  1489 => (x"26",x"87",x"d9",x"f9"),
  1490 => (x"0e",x"4f",x"26",x"4b"),
  1491 => (x"5d",x"5c",x"5b",x"5e"),
  1492 => (x"86",x"d4",x"ff",x"0e"),
  1493 => (x"c8",x"59",x"a6",x"dc"),
  1494 => (x"78",x"c0",x"48",x"a6"),
  1495 => (x"c0",x"c1",x"80",x"c4"),
  1496 => (x"80",x"c4",x"78",x"66"),
  1497 => (x"80",x"c4",x"78",x"c1"),
  1498 => (x"cd",x"c4",x"78",x"c1"),
  1499 => (x"78",x"c1",x"48",x"e8"),
  1500 => (x"bf",x"d8",x"cc",x"c4"),
  1501 => (x"05",x"a8",x"de",x"48"),
  1502 => (x"f6",x"f4",x"87",x"c9"),
  1503 => (x"58",x"a6",x"cc",x"87"),
  1504 => (x"c1",x"87",x"df",x"cf"),
  1505 => (x"e4",x"87",x"f4",x"f7"),
  1506 => (x"f7",x"c1",x"87",x"ec"),
  1507 => (x"4c",x"70",x"87",x"ca"),
  1508 => (x"02",x"ac",x"fb",x"c0"),
  1509 => (x"d8",x"87",x"f0",x"c1"),
  1510 => (x"e2",x"c1",x"05",x"66"),
  1511 => (x"66",x"fc",x"c0",x"87"),
  1512 => (x"6a",x"82",x"c4",x"4a"),
  1513 => (x"d8",x"ee",x"c1",x"7e"),
  1514 => (x"20",x"49",x"6e",x"48"),
  1515 => (x"10",x"41",x"20",x"41"),
  1516 => (x"66",x"fc",x"c0",x"51"),
  1517 => (x"c6",x"d8",x"c1",x"48"),
  1518 => (x"c7",x"49",x"6a",x"78"),
  1519 => (x"c0",x"51",x"74",x"81"),
  1520 => (x"c8",x"49",x"66",x"fc"),
  1521 => (x"c0",x"51",x"c1",x"81"),
  1522 => (x"c9",x"49",x"66",x"fc"),
  1523 => (x"c0",x"51",x"c0",x"81"),
  1524 => (x"ca",x"49",x"66",x"fc"),
  1525 => (x"c1",x"51",x"c0",x"81"),
  1526 => (x"6a",x"1e",x"d8",x"1e"),
  1527 => (x"e3",x"81",x"c8",x"49"),
  1528 => (x"86",x"c8",x"87",x"e9"),
  1529 => (x"48",x"66",x"c0",x"c1"),
  1530 => (x"c7",x"01",x"a8",x"c0"),
  1531 => (x"48",x"a6",x"c8",x"87"),
  1532 => (x"87",x"ce",x"78",x"c1"),
  1533 => (x"48",x"66",x"c0",x"c1"),
  1534 => (x"a6",x"d0",x"88",x"c1"),
  1535 => (x"e2",x"87",x"c3",x"58"),
  1536 => (x"a6",x"d0",x"87",x"f4"),
  1537 => (x"74",x"78",x"c2",x"48"),
  1538 => (x"d1",x"cd",x"02",x"9c"),
  1539 => (x"48",x"66",x"c8",x"87"),
  1540 => (x"a8",x"66",x"c4",x"c1"),
  1541 => (x"87",x"c6",x"cd",x"03"),
  1542 => (x"c0",x"48",x"a6",x"dc"),
  1543 => (x"f4",x"c1",x"7e",x"78"),
  1544 => (x"4c",x"70",x"87",x"f6"),
  1545 => (x"05",x"ac",x"d0",x"c1"),
  1546 => (x"c4",x"87",x"d9",x"c2"),
  1547 => (x"78",x"6e",x"48",x"a6"),
  1548 => (x"70",x"87",x"c5",x"e4"),
  1549 => (x"df",x"f4",x"c1",x"7e"),
  1550 => (x"c0",x"4c",x"70",x"87"),
  1551 => (x"c1",x"05",x"ac",x"ec"),
  1552 => (x"66",x"c8",x"87",x"ed"),
  1553 => (x"c0",x"91",x"cc",x"49"),
  1554 => (x"c4",x"81",x"66",x"fc"),
  1555 => (x"4d",x"6a",x"4a",x"a1"),
  1556 => (x"6e",x"4a",x"a1",x"c8"),
  1557 => (x"ec",x"d1",x"c1",x"52"),
  1558 => (x"fb",x"f3",x"c1",x"79"),
  1559 => (x"9c",x"4c",x"70",x"87"),
  1560 => (x"c0",x"87",x"d9",x"02"),
  1561 => (x"d3",x"02",x"ac",x"fb"),
  1562 => (x"c1",x"55",x"74",x"87"),
  1563 => (x"70",x"87",x"e9",x"f3"),
  1564 => (x"c7",x"02",x"9c",x"4c"),
  1565 => (x"ac",x"fb",x"c0",x"87"),
  1566 => (x"87",x"ed",x"ff",x"05"),
  1567 => (x"c2",x"55",x"e0",x"c0"),
  1568 => (x"97",x"c0",x"55",x"c1"),
  1569 => (x"48",x"66",x"d8",x"7d"),
  1570 => (x"05",x"a8",x"66",x"c4"),
  1571 => (x"66",x"c8",x"87",x"db"),
  1572 => (x"a8",x"66",x"cc",x"48"),
  1573 => (x"c8",x"87",x"ca",x"04"),
  1574 => (x"80",x"c1",x"48",x"66"),
  1575 => (x"c8",x"58",x"a6",x"cc"),
  1576 => (x"48",x"66",x"cc",x"87"),
  1577 => (x"a6",x"d0",x"88",x"c1"),
  1578 => (x"eb",x"f2",x"c1",x"58"),
  1579 => (x"c1",x"4c",x"70",x"87"),
  1580 => (x"c8",x"05",x"ac",x"d0"),
  1581 => (x"48",x"66",x"d4",x"87"),
  1582 => (x"a6",x"d8",x"80",x"c1"),
  1583 => (x"ac",x"d0",x"c1",x"58"),
  1584 => (x"87",x"e7",x"fd",x"02"),
  1585 => (x"66",x"d8",x"48",x"6e"),
  1586 => (x"e3",x"c9",x"05",x"a8"),
  1587 => (x"a6",x"e0",x"c0",x"87"),
  1588 => (x"74",x"78",x"c0",x"48"),
  1589 => (x"88",x"fb",x"c0",x"48"),
  1590 => (x"70",x"58",x"a6",x"c8"),
  1591 => (x"e4",x"c9",x"02",x"98"),
  1592 => (x"88",x"cb",x"48",x"87"),
  1593 => (x"70",x"58",x"a6",x"c8"),
  1594 => (x"d1",x"c1",x"02",x"98"),
  1595 => (x"88",x"c9",x"48",x"87"),
  1596 => (x"70",x"58",x"a6",x"c8"),
  1597 => (x"c1",x"c4",x"02",x"98"),
  1598 => (x"88",x"c4",x"48",x"87"),
  1599 => (x"70",x"58",x"a6",x"c8"),
  1600 => (x"87",x"cf",x"02",x"98"),
  1601 => (x"c8",x"88",x"c1",x"48"),
  1602 => (x"98",x"70",x"58",x"a6"),
  1603 => (x"87",x"ea",x"c3",x"02"),
  1604 => (x"dc",x"87",x"d4",x"c8"),
  1605 => (x"f0",x"c0",x"48",x"a6"),
  1606 => (x"fb",x"f0",x"c1",x"78"),
  1607 => (x"c0",x"4c",x"70",x"87"),
  1608 => (x"c0",x"02",x"ac",x"ec"),
  1609 => (x"e0",x"c0",x"87",x"c4"),
  1610 => (x"ec",x"c0",x"5c",x"a6"),
  1611 => (x"cd",x"c0",x"02",x"ac"),
  1612 => (x"e3",x"f0",x"c1",x"87"),
  1613 => (x"c0",x"4c",x"70",x"87"),
  1614 => (x"ff",x"05",x"ac",x"ec"),
  1615 => (x"ec",x"c0",x"87",x"f3"),
  1616 => (x"c4",x"c0",x"02",x"ac"),
  1617 => (x"cf",x"f0",x"c1",x"87"),
  1618 => (x"ca",x"1e",x"c0",x"87"),
  1619 => (x"49",x"66",x"d0",x"1e"),
  1620 => (x"c4",x"c1",x"91",x"cc"),
  1621 => (x"80",x"71",x"48",x"66"),
  1622 => (x"c8",x"58",x"a6",x"cc"),
  1623 => (x"80",x"c4",x"48",x"66"),
  1624 => (x"cc",x"58",x"a6",x"d0"),
  1625 => (x"ff",x"49",x"bf",x"66"),
  1626 => (x"c1",x"87",x"e0",x"dd"),
  1627 => (x"d4",x"1e",x"de",x"1e"),
  1628 => (x"ff",x"49",x"bf",x"66"),
  1629 => (x"d0",x"87",x"d4",x"dd"),
  1630 => (x"48",x"49",x"70",x"86"),
  1631 => (x"c0",x"88",x"08",x"c0"),
  1632 => (x"c0",x"58",x"a6",x"e8"),
  1633 => (x"ee",x"c0",x"06",x"a8"),
  1634 => (x"66",x"e4",x"c0",x"87"),
  1635 => (x"03",x"a8",x"dd",x"48"),
  1636 => (x"c4",x"87",x"e4",x"c0"),
  1637 => (x"c0",x"49",x"bf",x"66"),
  1638 => (x"c0",x"81",x"66",x"e4"),
  1639 => (x"e4",x"c0",x"51",x"e0"),
  1640 => (x"81",x"c1",x"49",x"66"),
  1641 => (x"81",x"bf",x"66",x"c4"),
  1642 => (x"c0",x"51",x"c1",x"c2"),
  1643 => (x"c2",x"49",x"66",x"e4"),
  1644 => (x"bf",x"66",x"c4",x"81"),
  1645 => (x"6e",x"51",x"c0",x"81"),
  1646 => (x"c6",x"d8",x"c1",x"48"),
  1647 => (x"c8",x"49",x"6e",x"78"),
  1648 => (x"51",x"66",x"d0",x"81"),
  1649 => (x"81",x"c9",x"49",x"6e"),
  1650 => (x"6e",x"51",x"66",x"d4"),
  1651 => (x"dc",x"81",x"ca",x"49"),
  1652 => (x"66",x"d0",x"51",x"66"),
  1653 => (x"d4",x"80",x"c1",x"48"),
  1654 => (x"66",x"c8",x"58",x"a6"),
  1655 => (x"a8",x"66",x"cc",x"48"),
  1656 => (x"87",x"cb",x"c0",x"04"),
  1657 => (x"c1",x"48",x"66",x"c8"),
  1658 => (x"58",x"a6",x"cc",x"80"),
  1659 => (x"cc",x"87",x"d6",x"c5"),
  1660 => (x"88",x"c1",x"48",x"66"),
  1661 => (x"c5",x"58",x"a6",x"d0"),
  1662 => (x"dc",x"ff",x"87",x"cb"),
  1663 => (x"e8",x"c0",x"87",x"fa"),
  1664 => (x"dc",x"ff",x"58",x"a6"),
  1665 => (x"e0",x"c0",x"87",x"f2"),
  1666 => (x"ec",x"c0",x"58",x"a6"),
  1667 => (x"ca",x"c0",x"05",x"a8"),
  1668 => (x"48",x"a6",x"dc",x"87"),
  1669 => (x"78",x"66",x"e4",x"c0"),
  1670 => (x"c1",x"87",x"c4",x"c0"),
  1671 => (x"c8",x"87",x"f9",x"ec"),
  1672 => (x"91",x"cc",x"49",x"66"),
  1673 => (x"48",x"66",x"fc",x"c0"),
  1674 => (x"a6",x"c8",x"80",x"71"),
  1675 => (x"4a",x"66",x"c4",x"58"),
  1676 => (x"66",x"c4",x"82",x"c8"),
  1677 => (x"c0",x"81",x"ca",x"49"),
  1678 => (x"dc",x"51",x"66",x"e4"),
  1679 => (x"81",x"c1",x"49",x"66"),
  1680 => (x"89",x"66",x"e4",x"c0"),
  1681 => (x"30",x"71",x"48",x"c1"),
  1682 => (x"89",x"c1",x"49",x"70"),
  1683 => (x"c4",x"7a",x"97",x"71"),
  1684 => (x"49",x"bf",x"f4",x"d1"),
  1685 => (x"29",x"66",x"e4",x"c0"),
  1686 => (x"48",x"4a",x"6a",x"97"),
  1687 => (x"ec",x"c0",x"98",x"71"),
  1688 => (x"66",x"c4",x"58",x"a6"),
  1689 => (x"69",x"81",x"c4",x"49"),
  1690 => (x"48",x"66",x"d8",x"4d"),
  1691 => (x"c0",x"02",x"a8",x"6e"),
  1692 => (x"7e",x"c0",x"87",x"c5"),
  1693 => (x"c1",x"87",x"c2",x"c0"),
  1694 => (x"c0",x"1e",x"6e",x"7e"),
  1695 => (x"49",x"75",x"1e",x"e0"),
  1696 => (x"87",x"c7",x"d9",x"ff"),
  1697 => (x"4c",x"70",x"86",x"c8"),
  1698 => (x"06",x"ac",x"b7",x"c0"),
  1699 => (x"74",x"87",x"d0",x"c1"),
  1700 => (x"49",x"e0",x"c0",x"85"),
  1701 => (x"4b",x"75",x"89",x"74"),
  1702 => (x"4a",x"e4",x"ee",x"c1"),
  1703 => (x"e1",x"d8",x"fe",x"71"),
  1704 => (x"75",x"85",x"c2",x"87"),
  1705 => (x"66",x"e0",x"c0",x"7e"),
  1706 => (x"c0",x"80",x"c1",x"48"),
  1707 => (x"c0",x"58",x"a6",x"e4"),
  1708 => (x"c1",x"49",x"66",x"e8"),
  1709 => (x"02",x"a9",x"70",x"81"),
  1710 => (x"c0",x"87",x"c5",x"c0"),
  1711 => (x"87",x"c2",x"c0",x"4d"),
  1712 => (x"1e",x"75",x"4d",x"c1"),
  1713 => (x"c0",x"49",x"a4",x"c2"),
  1714 => (x"88",x"71",x"48",x"e0"),
  1715 => (x"c8",x"1e",x"49",x"70"),
  1716 => (x"d7",x"ff",x"49",x"66"),
  1717 => (x"86",x"c8",x"87",x"f5"),
  1718 => (x"01",x"a8",x"b7",x"c0"),
  1719 => (x"c0",x"87",x"c6",x"ff"),
  1720 => (x"c0",x"02",x"66",x"e0"),
  1721 => (x"66",x"c4",x"87",x"d3"),
  1722 => (x"c0",x"81",x"c9",x"49"),
  1723 => (x"c4",x"51",x"66",x"e0"),
  1724 => (x"d9",x"c1",x"48",x"66"),
  1725 => (x"ce",x"c0",x"78",x"ca"),
  1726 => (x"49",x"66",x"c4",x"87"),
  1727 => (x"51",x"c2",x"81",x"c9"),
  1728 => (x"c3",x"48",x"66",x"c4"),
  1729 => (x"c8",x"78",x"d8",x"dd"),
  1730 => (x"66",x"cc",x"48",x"66"),
  1731 => (x"cb",x"c0",x"04",x"a8"),
  1732 => (x"48",x"66",x"c8",x"87"),
  1733 => (x"a6",x"cc",x"80",x"c1"),
  1734 => (x"87",x"e9",x"c0",x"58"),
  1735 => (x"c1",x"48",x"66",x"cc"),
  1736 => (x"58",x"a6",x"d0",x"88"),
  1737 => (x"ff",x"87",x"de",x"c0"),
  1738 => (x"70",x"87",x"cb",x"d6"),
  1739 => (x"87",x"d5",x"c0",x"4c"),
  1740 => (x"05",x"ac",x"c6",x"c1"),
  1741 => (x"d0",x"87",x"c8",x"c0"),
  1742 => (x"80",x"c1",x"48",x"66"),
  1743 => (x"ff",x"58",x"a6",x"d4"),
  1744 => (x"70",x"87",x"f3",x"d5"),
  1745 => (x"48",x"66",x"d4",x"4c"),
  1746 => (x"a6",x"d8",x"80",x"c1"),
  1747 => (x"02",x"9c",x"74",x"58"),
  1748 => (x"c8",x"87",x"cb",x"c0"),
  1749 => (x"c4",x"c1",x"48",x"66"),
  1750 => (x"f2",x"04",x"a8",x"66"),
  1751 => (x"d5",x"ff",x"87",x"fa"),
  1752 => (x"66",x"c8",x"87",x"cb"),
  1753 => (x"03",x"a8",x"c7",x"48"),
  1754 => (x"c8",x"87",x"e1",x"c0"),
  1755 => (x"cd",x"c4",x"4c",x"66"),
  1756 => (x"78",x"c0",x"48",x"e8"),
  1757 => (x"91",x"cc",x"49",x"74"),
  1758 => (x"81",x"66",x"fc",x"c0"),
  1759 => (x"6a",x"4a",x"a1",x"c4"),
  1760 => (x"79",x"52",x"c0",x"4a"),
  1761 => (x"ac",x"c7",x"84",x"c1"),
  1762 => (x"87",x"e2",x"ff",x"04"),
  1763 => (x"26",x"8e",x"d4",x"ff"),
  1764 => (x"26",x"4c",x"26",x"4d"),
  1765 => (x"00",x"4f",x"26",x"4b"),
  1766 => (x"64",x"61",x"6f",x"4c"),
  1767 => (x"20",x"2e",x"2a",x"20"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"1e",x"00",x"20",x"3a"),
  1770 => (x"4b",x"71",x"1e",x"73"),
  1771 => (x"87",x"c6",x"02",x"9b"),
  1772 => (x"48",x"e4",x"cd",x"c4"),
  1773 => (x"1e",x"c7",x"78",x"c0"),
  1774 => (x"bf",x"e4",x"cd",x"c4"),
  1775 => (x"fc",x"f3",x"c1",x"1e"),
  1776 => (x"d8",x"cc",x"c4",x"1e"),
  1777 => (x"c2",x"ee",x"49",x"bf"),
  1778 => (x"c4",x"86",x"cc",x"87"),
  1779 => (x"49",x"bf",x"d8",x"cc"),
  1780 => (x"73",x"87",x"f8",x"e2"),
  1781 => (x"87",x"c8",x"02",x"9b"),
  1782 => (x"49",x"fc",x"f3",x"c1"),
  1783 => (x"87",x"ce",x"e8",x"c0"),
  1784 => (x"4f",x"26",x"4b",x"26"),
  1785 => (x"fc",x"1e",x"73",x"1e"),
  1786 => (x"4b",x"ff",x"c3",x"86"),
  1787 => (x"fc",x"4a",x"d4",x"ff"),
  1788 => (x"98",x"c1",x"48",x"bf"),
  1789 => (x"98",x"48",x"7e",x"70"),
  1790 => (x"87",x"fb",x"c0",x"02"),
  1791 => (x"c1",x"48",x"d0",x"ff"),
  1792 => (x"d2",x"c2",x"78",x"c1"),
  1793 => (x"c3",x"7a",x"73",x"7a"),
  1794 => (x"48",x"49",x"e1",x"ff"),
  1795 => (x"50",x"6a",x"80",x"ff"),
  1796 => (x"51",x"6a",x"7a",x"73"),
  1797 => (x"80",x"c1",x"7a",x"73"),
  1798 => (x"7a",x"73",x"50",x"6a"),
  1799 => (x"7a",x"73",x"50",x"6a"),
  1800 => (x"7a",x"73",x"49",x"6a"),
  1801 => (x"7a",x"73",x"50",x"6a"),
  1802 => (x"ff",x"c3",x"50",x"6a"),
  1803 => (x"ff",x"59",x"97",x"ea"),
  1804 => (x"c0",x"c1",x"48",x"d0"),
  1805 => (x"c3",x"87",x"d7",x"78"),
  1806 => (x"48",x"49",x"e1",x"ff"),
  1807 => (x"50",x"c0",x"80",x"ff"),
  1808 => (x"c0",x"80",x"c1",x"51"),
  1809 => (x"c1",x"50",x"d9",x"50"),
  1810 => (x"50",x"e2",x"c0",x"50"),
  1811 => (x"ff",x"c3",x"50",x"c3"),
  1812 => (x"50",x"c0",x"48",x"e7"),
  1813 => (x"8e",x"fc",x"80",x"f8"),
  1814 => (x"4f",x"26",x"4b",x"26"),
  1815 => (x"87",x"d5",x"cc",x"1e"),
  1816 => (x"c2",x"fd",x"49",x"c1"),
  1817 => (x"d1",x"dc",x"fe",x"87"),
  1818 => (x"02",x"98",x"70",x"87"),
  1819 => (x"e5",x"fe",x"87",x"cd"),
  1820 => (x"98",x"70",x"87",x"dd"),
  1821 => (x"c1",x"87",x"c4",x"02"),
  1822 => (x"c0",x"87",x"c2",x"4a"),
  1823 => (x"05",x"9a",x"72",x"4a"),
  1824 => (x"1e",x"c0",x"87",x"ce"),
  1825 => (x"49",x"f0",x"f2",x"c1"),
  1826 => (x"87",x"ed",x"f2",x"c0"),
  1827 => (x"87",x"fe",x"86",x"c4"),
  1828 => (x"f2",x"c1",x"1e",x"c0"),
  1829 => (x"f2",x"c0",x"49",x"fc"),
  1830 => (x"1e",x"c0",x"87",x"df"),
  1831 => (x"87",x"d1",x"f9",x"c1"),
  1832 => (x"f2",x"c0",x"49",x"70"),
  1833 => (x"d7",x"c3",x"87",x"d3"),
  1834 => (x"26",x"8e",x"f8",x"87"),
  1835 => (x"00",x"00",x"00",x"4f"),
  1836 => (x"66",x"20",x"44",x"53"),
  1837 => (x"65",x"6c",x"69",x"61"),
  1838 => (x"00",x"00",x"2e",x"64"),
  1839 => (x"74",x"6f",x"6f",x"42"),
  1840 => (x"2e",x"67",x"6e",x"69"),
  1841 => (x"1e",x"00",x"2e",x"2e"),
  1842 => (x"48",x"e4",x"cd",x"c4"),
  1843 => (x"cc",x"c4",x"78",x"c0"),
  1844 => (x"78",x"c0",x"48",x"d8"),
  1845 => (x"c1",x"87",x"c5",x"fe"),
  1846 => (x"c0",x"87",x"f3",x"fb"),
  1847 => (x"00",x"4f",x"26",x"48"),
  1848 => (x"00",x"00",x"00",x"00"),
  1849 => (x"00",x"00",x"00",x"00"),
  1850 => (x"00",x"00",x"00",x"01"),
  1851 => (x"78",x"45",x"20",x"80"),
  1852 => (x"00",x"00",x"74",x"69"),
  1853 => (x"61",x"42",x"20",x"80"),
  1854 => (x"00",x"00",x"6b",x"63"),
  1855 => (x"00",x"00",x"13",x"ad"),
  1856 => (x"00",x"00",x"43",x"78"),
  1857 => (x"00",x"00",x"00",x"00"),
  1858 => (x"00",x"00",x"13",x"ad"),
  1859 => (x"00",x"00",x"43",x"96"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"13",x"ad"),
  1862 => (x"00",x"00",x"43",x"b4"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"13",x"ad"),
  1865 => (x"00",x"00",x"43",x"d2"),
  1866 => (x"00",x"00",x"00",x"00"),
  1867 => (x"00",x"00",x"13",x"ad"),
  1868 => (x"00",x"00",x"43",x"f0"),
  1869 => (x"00",x"00",x"00",x"00"),
  1870 => (x"00",x"00",x"13",x"ad"),
  1871 => (x"00",x"00",x"44",x"0e"),
  1872 => (x"00",x"00",x"00",x"00"),
  1873 => (x"00",x"00",x"13",x"ad"),
  1874 => (x"00",x"00",x"44",x"2c"),
  1875 => (x"00",x"00",x"00",x"00"),
  1876 => (x"00",x"00",x"14",x"6c"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"16",x"bb"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"48",x"f0",x"fe",x"1e"),
  1883 => (x"09",x"cd",x"78",x"c0"),
  1884 => (x"4f",x"26",x"09",x"79"),
  1885 => (x"fe",x"86",x"fc",x"1e"),
  1886 => (x"48",x"7e",x"bf",x"f0"),
  1887 => (x"4f",x"26",x"8e",x"fc"),
  1888 => (x"48",x"f0",x"fe",x"1e"),
  1889 => (x"4f",x"26",x"78",x"c1"),
  1890 => (x"48",x"f0",x"fe",x"1e"),
  1891 => (x"4f",x"26",x"78",x"c0"),
  1892 => (x"c0",x"4a",x"71",x"1e"),
  1893 => (x"a2",x"c1",x"7a",x"97"),
  1894 => (x"ca",x"51",x"c0",x"49"),
  1895 => (x"51",x"c0",x"49",x"a2"),
  1896 => (x"c0",x"49",x"a2",x"cb"),
  1897 => (x"0e",x"4f",x"26",x"51"),
  1898 => (x"0e",x"5c",x"5b",x"5e"),
  1899 => (x"4c",x"71",x"86",x"f0"),
  1900 => (x"97",x"49",x"a4",x"ca"),
  1901 => (x"a4",x"cb",x"7e",x"69"),
  1902 => (x"48",x"6b",x"97",x"4b"),
  1903 => (x"c1",x"58",x"a6",x"c8"),
  1904 => (x"58",x"a6",x"cc",x"80"),
  1905 => (x"a6",x"d0",x"98",x"c7"),
  1906 => (x"cc",x"48",x"6e",x"58"),
  1907 => (x"db",x"05",x"a8",x"66"),
  1908 => (x"7e",x"69",x"97",x"87"),
  1909 => (x"c8",x"48",x"6b",x"97"),
  1910 => (x"80",x"c1",x"58",x"a6"),
  1911 => (x"c7",x"58",x"a6",x"cc"),
  1912 => (x"58",x"a6",x"d0",x"98"),
  1913 => (x"66",x"cc",x"48",x"6e"),
  1914 => (x"87",x"e5",x"02",x"a8"),
  1915 => (x"cc",x"87",x"d9",x"fe"),
  1916 => (x"6b",x"97",x"4a",x"a4"),
  1917 => (x"49",x"a1",x"72",x"49"),
  1918 => (x"97",x"51",x"66",x"dc"),
  1919 => (x"48",x"6e",x"7e",x"6b"),
  1920 => (x"a6",x"c8",x"80",x"c1"),
  1921 => (x"cc",x"98",x"c7",x"58"),
  1922 => (x"97",x"70",x"58",x"a6"),
  1923 => (x"87",x"d1",x"c2",x"7b"),
  1924 => (x"f0",x"87",x"ed",x"fd"),
  1925 => (x"26",x"4c",x"26",x"8e"),
  1926 => (x"0e",x"4f",x"26",x"4b"),
  1927 => (x"5d",x"5c",x"5b",x"5e"),
  1928 => (x"71",x"86",x"f4",x"0e"),
  1929 => (x"7e",x"6d",x"97",x"4d"),
  1930 => (x"97",x"4c",x"a5",x"c1"),
  1931 => (x"a6",x"c8",x"48",x"6c"),
  1932 => (x"c4",x"48",x"6e",x"58"),
  1933 => (x"c5",x"05",x"a8",x"66"),
  1934 => (x"c0",x"48",x"ff",x"87"),
  1935 => (x"c7",x"fd",x"87",x"e6"),
  1936 => (x"49",x"a5",x"c2",x"87"),
  1937 => (x"71",x"4b",x"6c",x"97"),
  1938 => (x"6b",x"97",x"4b",x"a3"),
  1939 => (x"7e",x"6c",x"97",x"4b"),
  1940 => (x"80",x"c1",x"48",x"6e"),
  1941 => (x"c7",x"58",x"a6",x"c8"),
  1942 => (x"58",x"a6",x"cc",x"98"),
  1943 => (x"fc",x"7c",x"97",x"70"),
  1944 => (x"48",x"73",x"87",x"de"),
  1945 => (x"4d",x"26",x"8e",x"f4"),
  1946 => (x"4b",x"26",x"4c",x"26"),
  1947 => (x"5e",x"0e",x"4f",x"26"),
  1948 => (x"f4",x"0e",x"5c",x"5b"),
  1949 => (x"d8",x"4c",x"71",x"86"),
  1950 => (x"ff",x"c3",x"4a",x"66"),
  1951 => (x"4b",x"a4",x"c2",x"9a"),
  1952 => (x"73",x"49",x"6c",x"97"),
  1953 => (x"51",x"72",x"49",x"a1"),
  1954 => (x"6e",x"7e",x"6c",x"97"),
  1955 => (x"c8",x"80",x"c1",x"48"),
  1956 => (x"98",x"c7",x"58",x"a6"),
  1957 => (x"70",x"58",x"a6",x"cc"),
  1958 => (x"26",x"8e",x"f4",x"54"),
  1959 => (x"26",x"4b",x"26",x"4c"),
  1960 => (x"1e",x"73",x"1e",x"4f"),
  1961 => (x"df",x"fb",x"86",x"f4"),
  1962 => (x"4b",x"bf",x"e0",x"87"),
  1963 => (x"c0",x"e0",x"c0",x"49"),
  1964 => (x"87",x"cb",x"02",x"99"),
  1965 => (x"d1",x"c4",x"1e",x"73"),
  1966 => (x"f1",x"fe",x"49",x"cc"),
  1967 => (x"73",x"86",x"c4",x"87"),
  1968 => (x"99",x"c0",x"d0",x"49"),
  1969 => (x"87",x"c0",x"c1",x"02"),
  1970 => (x"97",x"d6",x"d1",x"c4"),
  1971 => (x"d1",x"c4",x"7e",x"bf"),
  1972 => (x"48",x"bf",x"97",x"d7"),
  1973 => (x"6e",x"58",x"a6",x"c8"),
  1974 => (x"a8",x"66",x"c4",x"48"),
  1975 => (x"87",x"e8",x"c0",x"02"),
  1976 => (x"97",x"d6",x"d1",x"c4"),
  1977 => (x"d1",x"c4",x"49",x"bf"),
  1978 => (x"48",x"11",x"81",x"d8"),
  1979 => (x"c4",x"78",x"08",x"e0"),
  1980 => (x"bf",x"97",x"d6",x"d1"),
  1981 => (x"c1",x"48",x"6e",x"7e"),
  1982 => (x"58",x"a6",x"c8",x"80"),
  1983 => (x"a6",x"cc",x"98",x"c7"),
  1984 => (x"d6",x"d1",x"c4",x"58"),
  1985 => (x"50",x"66",x"c8",x"48"),
  1986 => (x"49",x"4b",x"bf",x"e4"),
  1987 => (x"99",x"c0",x"e0",x"c0"),
  1988 => (x"73",x"87",x"cb",x"02"),
  1989 => (x"e0",x"d1",x"c4",x"1e"),
  1990 => (x"87",x"d2",x"fd",x"49"),
  1991 => (x"49",x"73",x"86",x"c4"),
  1992 => (x"02",x"99",x"c0",x"d0"),
  1993 => (x"c4",x"87",x"c0",x"c1"),
  1994 => (x"bf",x"97",x"ea",x"d1"),
  1995 => (x"eb",x"d1",x"c4",x"7e"),
  1996 => (x"c8",x"48",x"bf",x"97"),
  1997 => (x"48",x"6e",x"58",x"a6"),
  1998 => (x"02",x"a8",x"66",x"c4"),
  1999 => (x"c4",x"87",x"e8",x"c0"),
  2000 => (x"bf",x"97",x"ea",x"d1"),
  2001 => (x"ec",x"d1",x"c4",x"49"),
  2002 => (x"e4",x"48",x"11",x"81"),
  2003 => (x"d1",x"c4",x"78",x"08"),
  2004 => (x"7e",x"bf",x"97",x"ea"),
  2005 => (x"80",x"c1",x"48",x"6e"),
  2006 => (x"c7",x"58",x"a6",x"c8"),
  2007 => (x"58",x"a6",x"cc",x"98"),
  2008 => (x"48",x"ea",x"d1",x"c4"),
  2009 => (x"f8",x"50",x"66",x"c8"),
  2010 => (x"7e",x"70",x"87",x"ca"),
  2011 => (x"f4",x"87",x"d1",x"f8"),
  2012 => (x"26",x"4b",x"26",x"8e"),
  2013 => (x"d1",x"c4",x"1e",x"4f"),
  2014 => (x"d3",x"f8",x"49",x"cc"),
  2015 => (x"e0",x"d1",x"c4",x"87"),
  2016 => (x"87",x"cc",x"f8",x"49"),
  2017 => (x"49",x"e1",x"fa",x"c1"),
  2018 => (x"c2",x"87",x"dd",x"f7"),
  2019 => (x"4f",x"26",x"87",x"f2"),
  2020 => (x"c4",x"1e",x"73",x"1e"),
  2021 => (x"fa",x"49",x"cc",x"d1"),
  2022 => (x"4a",x"70",x"87",x"c1"),
  2023 => (x"04",x"aa",x"b7",x"c0"),
  2024 => (x"c3",x"87",x"cc",x"c2"),
  2025 => (x"c9",x"05",x"aa",x"f0"),
  2026 => (x"f8",x"c0",x"c2",x"87"),
  2027 => (x"c1",x"78",x"c1",x"48"),
  2028 => (x"e0",x"c3",x"87",x"ed"),
  2029 => (x"87",x"c9",x"05",x"aa"),
  2030 => (x"48",x"fc",x"c0",x"c2"),
  2031 => (x"de",x"c1",x"78",x"c1"),
  2032 => (x"fc",x"c0",x"c2",x"87"),
  2033 => (x"87",x"c6",x"02",x"bf"),
  2034 => (x"4b",x"a2",x"c0",x"c2"),
  2035 => (x"4b",x"72",x"87",x"c2"),
  2036 => (x"bf",x"f8",x"c0",x"c2"),
  2037 => (x"87",x"e0",x"c0",x"02"),
  2038 => (x"b7",x"c4",x"49",x"73"),
  2039 => (x"c2",x"c2",x"91",x"29"),
  2040 => (x"4a",x"73",x"81",x"d4"),
  2041 => (x"92",x"c2",x"9a",x"cf"),
  2042 => (x"30",x"72",x"48",x"c1"),
  2043 => (x"ba",x"ff",x"4a",x"70"),
  2044 => (x"98",x"69",x"48",x"72"),
  2045 => (x"87",x"db",x"79",x"70"),
  2046 => (x"b7",x"c4",x"49",x"73"),
  2047 => (x"c2",x"c2",x"91",x"29"),
  2048 => (x"4a",x"73",x"81",x"d4"),
  2049 => (x"92",x"c2",x"9a",x"cf"),
  2050 => (x"30",x"72",x"48",x"c3"),
  2051 => (x"69",x"48",x"4a",x"70"),
  2052 => (x"c2",x"79",x"70",x"b0"),
  2053 => (x"c0",x"48",x"fc",x"c0"),
  2054 => (x"f8",x"c0",x"c2",x"78"),
  2055 => (x"c4",x"78",x"c0",x"48"),
  2056 => (x"f7",x"49",x"cc",x"d1"),
  2057 => (x"4a",x"70",x"87",x"f5"),
  2058 => (x"03",x"aa",x"b7",x"c0"),
  2059 => (x"c0",x"87",x"f4",x"fd"),
  2060 => (x"26",x"4b",x"26",x"48"),
  2061 => (x"00",x"00",x"00",x"4f"),
  2062 => (x"00",x"00",x"00",x"00"),
  2063 => (x"00",x"00",x"00",x"00"),
  2064 => (x"72",x"4a",x"c0",x"1e"),
  2065 => (x"c2",x"91",x"c4",x"49"),
  2066 => (x"c0",x"81",x"d4",x"c2"),
  2067 => (x"d0",x"82",x"c1",x"79"),
  2068 => (x"ee",x"04",x"aa",x"b7"),
  2069 => (x"0e",x"4f",x"26",x"87"),
  2070 => (x"5d",x"5c",x"5b",x"5e"),
  2071 => (x"f4",x"4d",x"71",x"0e"),
  2072 => (x"4a",x"75",x"87",x"e6"),
  2073 => (x"92",x"2a",x"b7",x"c4"),
  2074 => (x"82",x"d4",x"c2",x"c2"),
  2075 => (x"9c",x"cf",x"4c",x"75"),
  2076 => (x"49",x"6a",x"94",x"c2"),
  2077 => (x"c3",x"2b",x"74",x"4b"),
  2078 => (x"74",x"48",x"c2",x"9b"),
  2079 => (x"ff",x"4c",x"70",x"30"),
  2080 => (x"71",x"48",x"74",x"bc"),
  2081 => (x"f3",x"7a",x"70",x"98"),
  2082 => (x"48",x"73",x"87",x"f6"),
  2083 => (x"4c",x"26",x"4d",x"26"),
  2084 => (x"4f",x"26",x"4b",x"26"),
  2085 => (x"00",x"00",x"00",x"00"),
  2086 => (x"00",x"00",x"00",x"00"),
  2087 => (x"00",x"00",x"00",x"00"),
  2088 => (x"00",x"00",x"00",x"00"),
  2089 => (x"00",x"00",x"00",x"00"),
  2090 => (x"00",x"00",x"00",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"00",x"00",x"00",x"00"),
  2093 => (x"00",x"00",x"00",x"00"),
  2094 => (x"00",x"00",x"00",x"00"),
  2095 => (x"00",x"00",x"00",x"00"),
  2096 => (x"00",x"00",x"00",x"00"),
  2097 => (x"00",x"00",x"00",x"00"),
  2098 => (x"00",x"00",x"00",x"00"),
  2099 => (x"00",x"00",x"00",x"00"),
  2100 => (x"00",x"00",x"00",x"00"),
  2101 => (x"48",x"d0",x"ff",x"1e"),
  2102 => (x"71",x"78",x"e1",x"c8"),
  2103 => (x"08",x"d4",x"ff",x"48"),
  2104 => (x"1e",x"4f",x"26",x"78"),
  2105 => (x"c8",x"48",x"d0",x"ff"),
  2106 => (x"48",x"71",x"78",x"e1"),
  2107 => (x"78",x"08",x"d4",x"ff"),
  2108 => (x"ff",x"48",x"66",x"c4"),
  2109 => (x"26",x"78",x"08",x"d4"),
  2110 => (x"4a",x"71",x"1e",x"4f"),
  2111 => (x"1e",x"49",x"66",x"c4"),
  2112 => (x"de",x"ff",x"49",x"72"),
  2113 => (x"48",x"d0",x"ff",x"87"),
  2114 => (x"fc",x"78",x"e0",x"c0"),
  2115 => (x"1e",x"4f",x"26",x"8e"),
  2116 => (x"4b",x"71",x"1e",x"73"),
  2117 => (x"1e",x"49",x"66",x"c8"),
  2118 => (x"e0",x"c1",x"4a",x"73"),
  2119 => (x"d8",x"ff",x"49",x"a2"),
  2120 => (x"26",x"8e",x"fc",x"87"),
  2121 => (x"1e",x"4f",x"26",x"4b"),
  2122 => (x"4b",x"71",x"1e",x"73"),
  2123 => (x"fe",x"49",x"e2",x"c0"),
  2124 => (x"4a",x"c7",x"87",x"e2"),
  2125 => (x"d4",x"ff",x"48",x"13"),
  2126 => (x"49",x"72",x"78",x"08"),
  2127 => (x"99",x"71",x"8a",x"c1"),
  2128 => (x"ff",x"87",x"f1",x"05"),
  2129 => (x"e0",x"c0",x"48",x"d0"),
  2130 => (x"26",x"4b",x"26",x"78"),
  2131 => (x"d0",x"ff",x"1e",x"4f"),
  2132 => (x"78",x"c9",x"c8",x"48"),
  2133 => (x"d4",x"ff",x"48",x"71"),
  2134 => (x"4f",x"26",x"78",x"08"),
  2135 => (x"49",x"4a",x"71",x"1e"),
  2136 => (x"d0",x"ff",x"87",x"eb"),
  2137 => (x"26",x"78",x"c8",x"48"),
  2138 => (x"1e",x"73",x"1e",x"4f"),
  2139 => (x"d2",x"c4",x"4b",x"71"),
  2140 => (x"c3",x"02",x"bf",x"c4"),
  2141 => (x"87",x"eb",x"c2",x"87"),
  2142 => (x"c8",x"48",x"d0",x"ff"),
  2143 => (x"48",x"73",x"78",x"c9"),
  2144 => (x"ff",x"b0",x"e0",x"c0"),
  2145 => (x"c4",x"78",x"08",x"d4"),
  2146 => (x"c0",x"48",x"f8",x"d1"),
  2147 => (x"02",x"66",x"c8",x"78"),
  2148 => (x"ff",x"c3",x"87",x"c5"),
  2149 => (x"c0",x"87",x"c2",x"49"),
  2150 => (x"c0",x"d2",x"c4",x"49"),
  2151 => (x"02",x"66",x"cc",x"59"),
  2152 => (x"d5",x"c5",x"87",x"c6"),
  2153 => (x"87",x"c4",x"4a",x"d5"),
  2154 => (x"4a",x"ff",x"ff",x"cf"),
  2155 => (x"5a",x"c4",x"d2",x"c4"),
  2156 => (x"48",x"c4",x"d2",x"c4"),
  2157 => (x"4b",x"26",x"78",x"c1"),
  2158 => (x"5e",x"0e",x"4f",x"26"),
  2159 => (x"0e",x"5d",x"5c",x"5b"),
  2160 => (x"d2",x"c4",x"4d",x"71"),
  2161 => (x"75",x"4b",x"bf",x"c0"),
  2162 => (x"87",x"cb",x"02",x"9d"),
  2163 => (x"c2",x"91",x"c8",x"49"),
  2164 => (x"71",x"4a",x"e0",x"c5"),
  2165 => (x"c2",x"87",x"c4",x"82"),
  2166 => (x"c0",x"4a",x"e0",x"c9"),
  2167 => (x"73",x"49",x"12",x"4c"),
  2168 => (x"fc",x"d1",x"c4",x"99"),
  2169 => (x"b8",x"71",x"48",x"bf"),
  2170 => (x"78",x"08",x"d4",x"ff"),
  2171 => (x"84",x"2b",x"b7",x"c1"),
  2172 => (x"04",x"ac",x"b7",x"c8"),
  2173 => (x"d1",x"c4",x"87",x"e7"),
  2174 => (x"c8",x"48",x"bf",x"f8"),
  2175 => (x"fc",x"d1",x"c4",x"80"),
  2176 => (x"26",x"4d",x"26",x"58"),
  2177 => (x"26",x"4b",x"26",x"4c"),
  2178 => (x"1e",x"73",x"1e",x"4f"),
  2179 => (x"4a",x"13",x"4b",x"71"),
  2180 => (x"87",x"cb",x"02",x"9a"),
  2181 => (x"e1",x"fe",x"49",x"72"),
  2182 => (x"9a",x"4a",x"13",x"87"),
  2183 => (x"26",x"87",x"f5",x"05"),
  2184 => (x"1e",x"4f",x"26",x"4b"),
  2185 => (x"bf",x"f8",x"d1",x"c4"),
  2186 => (x"f8",x"d1",x"c4",x"49"),
  2187 => (x"78",x"a1",x"c1",x"48"),
  2188 => (x"a9",x"b7",x"c0",x"c4"),
  2189 => (x"ff",x"87",x"db",x"03"),
  2190 => (x"d1",x"c4",x"48",x"d4"),
  2191 => (x"c4",x"78",x"bf",x"fc"),
  2192 => (x"49",x"bf",x"f8",x"d1"),
  2193 => (x"48",x"f8",x"d1",x"c4"),
  2194 => (x"c4",x"78",x"a1",x"c1"),
  2195 => (x"04",x"a9",x"b7",x"c0"),
  2196 => (x"d0",x"ff",x"87",x"e5"),
  2197 => (x"c4",x"78",x"c8",x"48"),
  2198 => (x"c0",x"48",x"c4",x"d2"),
  2199 => (x"00",x"4f",x"26",x"78"),
  2200 => (x"00",x"00",x"00",x"00"),
  2201 => (x"00",x"00",x"00",x"00"),
  2202 => (x"5f",x"00",x"00",x"00"),
  2203 => (x"00",x"00",x"00",x"5f"),
  2204 => (x"00",x"03",x"03",x"00"),
  2205 => (x"00",x"00",x"03",x"03"),
  2206 => (x"14",x"7f",x"7f",x"14"),
  2207 => (x"00",x"14",x"7f",x"7f"),
  2208 => (x"6b",x"2e",x"24",x"00"),
  2209 => (x"00",x"12",x"3a",x"6b"),
  2210 => (x"18",x"36",x"6a",x"4c"),
  2211 => (x"00",x"32",x"56",x"6c"),
  2212 => (x"59",x"4f",x"7e",x"30"),
  2213 => (x"40",x"68",x"3a",x"77"),
  2214 => (x"07",x"04",x"00",x"00"),
  2215 => (x"00",x"00",x"00",x"03"),
  2216 => (x"3e",x"1c",x"00",x"00"),
  2217 => (x"00",x"00",x"41",x"63"),
  2218 => (x"63",x"41",x"00",x"00"),
  2219 => (x"00",x"00",x"1c",x"3e"),
  2220 => (x"1c",x"3e",x"2a",x"08"),
  2221 => (x"08",x"2a",x"3e",x"1c"),
  2222 => (x"3e",x"08",x"08",x"00"),
  2223 => (x"00",x"08",x"08",x"3e"),
  2224 => (x"e0",x"80",x"00",x"00"),
  2225 => (x"00",x"00",x"00",x"60"),
  2226 => (x"08",x"08",x"08",x"00"),
  2227 => (x"00",x"08",x"08",x"08"),
  2228 => (x"60",x"00",x"00",x"00"),
  2229 => (x"00",x"00",x"00",x"60"),
  2230 => (x"18",x"30",x"60",x"40"),
  2231 => (x"01",x"03",x"06",x"0c"),
  2232 => (x"59",x"7f",x"3e",x"00"),
  2233 => (x"00",x"3e",x"7f",x"4d"),
  2234 => (x"7f",x"06",x"04",x"00"),
  2235 => (x"00",x"00",x"00",x"7f"),
  2236 => (x"71",x"63",x"42",x"00"),
  2237 => (x"00",x"46",x"4f",x"59"),
  2238 => (x"49",x"63",x"22",x"00"),
  2239 => (x"00",x"36",x"7f",x"49"),
  2240 => (x"13",x"16",x"1c",x"18"),
  2241 => (x"00",x"10",x"7f",x"7f"),
  2242 => (x"45",x"67",x"27",x"00"),
  2243 => (x"00",x"39",x"7d",x"45"),
  2244 => (x"4b",x"7e",x"3c",x"00"),
  2245 => (x"00",x"30",x"79",x"49"),
  2246 => (x"71",x"01",x"01",x"00"),
  2247 => (x"00",x"07",x"0f",x"79"),
  2248 => (x"49",x"7f",x"36",x"00"),
  2249 => (x"00",x"36",x"7f",x"49"),
  2250 => (x"49",x"4f",x"06",x"00"),
  2251 => (x"00",x"1e",x"3f",x"69"),
  2252 => (x"66",x"00",x"00",x"00"),
  2253 => (x"00",x"00",x"00",x"66"),
  2254 => (x"e6",x"80",x"00",x"00"),
  2255 => (x"00",x"00",x"00",x"66"),
  2256 => (x"14",x"08",x"08",x"00"),
  2257 => (x"00",x"22",x"22",x"14"),
  2258 => (x"14",x"14",x"14",x"00"),
  2259 => (x"00",x"14",x"14",x"14"),
  2260 => (x"14",x"22",x"22",x"00"),
  2261 => (x"00",x"08",x"08",x"14"),
  2262 => (x"51",x"03",x"02",x"00"),
  2263 => (x"00",x"06",x"0f",x"59"),
  2264 => (x"5d",x"41",x"7f",x"3e"),
  2265 => (x"00",x"1e",x"1f",x"55"),
  2266 => (x"09",x"7f",x"7e",x"00"),
  2267 => (x"00",x"7e",x"7f",x"09"),
  2268 => (x"49",x"7f",x"7f",x"00"),
  2269 => (x"00",x"36",x"7f",x"49"),
  2270 => (x"63",x"3e",x"1c",x"00"),
  2271 => (x"00",x"41",x"41",x"41"),
  2272 => (x"41",x"7f",x"7f",x"00"),
  2273 => (x"00",x"1c",x"3e",x"63"),
  2274 => (x"49",x"7f",x"7f",x"00"),
  2275 => (x"00",x"41",x"41",x"49"),
  2276 => (x"09",x"7f",x"7f",x"00"),
  2277 => (x"00",x"01",x"01",x"09"),
  2278 => (x"41",x"7f",x"3e",x"00"),
  2279 => (x"00",x"7a",x"7b",x"49"),
  2280 => (x"08",x"7f",x"7f",x"00"),
  2281 => (x"00",x"7f",x"7f",x"08"),
  2282 => (x"7f",x"41",x"00",x"00"),
  2283 => (x"00",x"00",x"41",x"7f"),
  2284 => (x"40",x"60",x"20",x"00"),
  2285 => (x"00",x"3f",x"7f",x"40"),
  2286 => (x"1c",x"08",x"7f",x"7f"),
  2287 => (x"00",x"41",x"63",x"36"),
  2288 => (x"40",x"7f",x"7f",x"00"),
  2289 => (x"00",x"40",x"40",x"40"),
  2290 => (x"0c",x"06",x"7f",x"7f"),
  2291 => (x"00",x"7f",x"7f",x"06"),
  2292 => (x"0c",x"06",x"7f",x"7f"),
  2293 => (x"00",x"7f",x"7f",x"18"),
  2294 => (x"41",x"7f",x"3e",x"00"),
  2295 => (x"00",x"3e",x"7f",x"41"),
  2296 => (x"09",x"7f",x"7f",x"00"),
  2297 => (x"00",x"06",x"0f",x"09"),
  2298 => (x"61",x"41",x"7f",x"3e"),
  2299 => (x"00",x"40",x"7e",x"7f"),
  2300 => (x"09",x"7f",x"7f",x"00"),
  2301 => (x"00",x"66",x"7f",x"19"),
  2302 => (x"4d",x"6f",x"26",x"00"),
  2303 => (x"00",x"32",x"7b",x"59"),
  2304 => (x"7f",x"01",x"01",x"00"),
  2305 => (x"00",x"01",x"01",x"7f"),
  2306 => (x"40",x"7f",x"3f",x"00"),
  2307 => (x"00",x"3f",x"7f",x"40"),
  2308 => (x"70",x"3f",x"0f",x"00"),
  2309 => (x"00",x"0f",x"3f",x"70"),
  2310 => (x"18",x"30",x"7f",x"7f"),
  2311 => (x"00",x"7f",x"7f",x"30"),
  2312 => (x"1c",x"36",x"63",x"41"),
  2313 => (x"41",x"63",x"36",x"1c"),
  2314 => (x"7c",x"06",x"03",x"01"),
  2315 => (x"01",x"03",x"06",x"7c"),
  2316 => (x"4d",x"59",x"71",x"61"),
  2317 => (x"00",x"41",x"43",x"47"),
  2318 => (x"7f",x"7f",x"00",x"00"),
  2319 => (x"00",x"00",x"41",x"41"),
  2320 => (x"0c",x"06",x"03",x"01"),
  2321 => (x"40",x"60",x"30",x"18"),
  2322 => (x"41",x"41",x"00",x"00"),
  2323 => (x"00",x"00",x"7f",x"7f"),
  2324 => (x"03",x"06",x"0c",x"08"),
  2325 => (x"00",x"08",x"0c",x"06"),
  2326 => (x"80",x"80",x"80",x"80"),
  2327 => (x"00",x"80",x"80",x"80"),
  2328 => (x"03",x"00",x"00",x"00"),
  2329 => (x"00",x"00",x"04",x"07"),
  2330 => (x"54",x"74",x"20",x"00"),
  2331 => (x"00",x"78",x"7c",x"54"),
  2332 => (x"44",x"7f",x"7f",x"00"),
  2333 => (x"00",x"38",x"7c",x"44"),
  2334 => (x"44",x"7c",x"38",x"00"),
  2335 => (x"00",x"00",x"44",x"44"),
  2336 => (x"44",x"7c",x"38",x"00"),
  2337 => (x"00",x"7f",x"7f",x"44"),
  2338 => (x"54",x"7c",x"38",x"00"),
  2339 => (x"00",x"18",x"5c",x"54"),
  2340 => (x"7f",x"7e",x"04",x"00"),
  2341 => (x"00",x"00",x"05",x"05"),
  2342 => (x"a4",x"bc",x"18",x"00"),
  2343 => (x"00",x"7c",x"fc",x"a4"),
  2344 => (x"04",x"7f",x"7f",x"00"),
  2345 => (x"00",x"78",x"7c",x"04"),
  2346 => (x"3d",x"00",x"00",x"00"),
  2347 => (x"00",x"00",x"40",x"7d"),
  2348 => (x"80",x"80",x"80",x"00"),
  2349 => (x"00",x"00",x"7d",x"fd"),
  2350 => (x"10",x"7f",x"7f",x"00"),
  2351 => (x"00",x"44",x"6c",x"38"),
  2352 => (x"3f",x"00",x"00",x"00"),
  2353 => (x"00",x"00",x"40",x"7f"),
  2354 => (x"18",x"0c",x"7c",x"7c"),
  2355 => (x"00",x"78",x"7c",x"0c"),
  2356 => (x"04",x"7c",x"7c",x"00"),
  2357 => (x"00",x"78",x"7c",x"04"),
  2358 => (x"44",x"7c",x"38",x"00"),
  2359 => (x"00",x"38",x"7c",x"44"),
  2360 => (x"24",x"fc",x"fc",x"00"),
  2361 => (x"00",x"18",x"3c",x"24"),
  2362 => (x"24",x"3c",x"18",x"00"),
  2363 => (x"00",x"fc",x"fc",x"24"),
  2364 => (x"04",x"7c",x"7c",x"00"),
  2365 => (x"00",x"08",x"0c",x"04"),
  2366 => (x"54",x"5c",x"48",x"00"),
  2367 => (x"00",x"20",x"74",x"54"),
  2368 => (x"7f",x"3f",x"04",x"00"),
  2369 => (x"00",x"00",x"44",x"44"),
  2370 => (x"40",x"7c",x"3c",x"00"),
  2371 => (x"00",x"7c",x"7c",x"40"),
  2372 => (x"60",x"3c",x"1c",x"00"),
  2373 => (x"00",x"1c",x"3c",x"60"),
  2374 => (x"30",x"60",x"7c",x"3c"),
  2375 => (x"00",x"3c",x"7c",x"60"),
  2376 => (x"10",x"38",x"6c",x"44"),
  2377 => (x"00",x"44",x"6c",x"38"),
  2378 => (x"e0",x"bc",x"1c",x"00"),
  2379 => (x"00",x"1c",x"3c",x"60"),
  2380 => (x"74",x"64",x"44",x"00"),
  2381 => (x"00",x"44",x"4c",x"5c"),
  2382 => (x"3e",x"08",x"08",x"00"),
  2383 => (x"00",x"41",x"41",x"77"),
  2384 => (x"7f",x"00",x"00",x"00"),
  2385 => (x"00",x"00",x"00",x"7f"),
  2386 => (x"77",x"41",x"41",x"00"),
  2387 => (x"00",x"08",x"08",x"3e"),
  2388 => (x"03",x"01",x"01",x"02"),
  2389 => (x"00",x"01",x"02",x"02"),
  2390 => (x"7f",x"7f",x"7f",x"7f"),
  2391 => (x"00",x"7f",x"7f",x"7f"),
  2392 => (x"1c",x"1c",x"08",x"08"),
  2393 => (x"7f",x"7f",x"3e",x"3e"),
  2394 => (x"3e",x"3e",x"7f",x"7f"),
  2395 => (x"08",x"08",x"1c",x"1c"),
  2396 => (x"7c",x"18",x"10",x"00"),
  2397 => (x"00",x"10",x"18",x"7c"),
  2398 => (x"7c",x"30",x"10",x"00"),
  2399 => (x"00",x"10",x"30",x"7c"),
  2400 => (x"60",x"60",x"30",x"10"),
  2401 => (x"00",x"06",x"1e",x"78"),
  2402 => (x"18",x"3c",x"66",x"42"),
  2403 => (x"00",x"42",x"66",x"3c"),
  2404 => (x"c2",x"6a",x"38",x"78"),
  2405 => (x"00",x"38",x"6c",x"c6"),
  2406 => (x"60",x"00",x"00",x"60"),
  2407 => (x"00",x"60",x"00",x"00"),
  2408 => (x"5c",x"5b",x"5e",x"0e"),
  2409 => (x"86",x"fc",x"0e",x"5d"),
  2410 => (x"d2",x"c4",x"7e",x"71"),
  2411 => (x"c0",x"4c",x"bf",x"d8"),
  2412 => (x"c4",x"1e",x"c0",x"4b"),
  2413 => (x"c4",x"02",x"ab",x"66"),
  2414 => (x"c2",x"4d",x"c0",x"87"),
  2415 => (x"75",x"4d",x"c1",x"87"),
  2416 => (x"ee",x"49",x"73",x"1e"),
  2417 => (x"86",x"c8",x"87",x"e3"),
  2418 => (x"ef",x"49",x"e0",x"c0"),
  2419 => (x"a4",x"c4",x"87",x"ec"),
  2420 => (x"f0",x"49",x"6a",x"4a"),
  2421 => (x"ca",x"f1",x"87",x"f3"),
  2422 => (x"c1",x"84",x"cc",x"87"),
  2423 => (x"ab",x"b7",x"c8",x"83"),
  2424 => (x"87",x"cd",x"ff",x"04"),
  2425 => (x"4d",x"26",x"8e",x"fc"),
  2426 => (x"4b",x"26",x"4c",x"26"),
  2427 => (x"71",x"1e",x"4f",x"26"),
  2428 => (x"dc",x"d2",x"c4",x"4a"),
  2429 => (x"dc",x"d2",x"c4",x"5a"),
  2430 => (x"49",x"78",x"c7",x"48"),
  2431 => (x"26",x"87",x"e1",x"fe"),
  2432 => (x"1e",x"73",x"1e",x"4f"),
  2433 => (x"b7",x"c0",x"4a",x"71"),
  2434 => (x"87",x"d3",x"03",x"aa"),
  2435 => (x"bf",x"dc",x"e6",x"c2"),
  2436 => (x"c1",x"87",x"c4",x"05"),
  2437 => (x"c0",x"87",x"c2",x"4b"),
  2438 => (x"e0",x"e6",x"c2",x"4b"),
  2439 => (x"c2",x"87",x"c4",x"5b"),
  2440 => (x"c2",x"5a",x"e0",x"e6"),
  2441 => (x"4a",x"bf",x"dc",x"e6"),
  2442 => (x"c0",x"c1",x"9a",x"c1"),
  2443 => (x"eb",x"ec",x"49",x"a2"),
  2444 => (x"c2",x"48",x"fc",x"87"),
  2445 => (x"78",x"bf",x"dc",x"e6"),
  2446 => (x"4f",x"26",x"4b",x"26"),
  2447 => (x"dc",x"e6",x"c2",x"1e"),
  2448 => (x"4f",x"26",x"48",x"bf"),
  2449 => (x"c4",x"4a",x"71",x"1e"),
  2450 => (x"49",x"72",x"1e",x"66"),
  2451 => (x"fc",x"87",x"c0",x"eb"),
  2452 => (x"1e",x"4f",x"26",x"8e"),
  2453 => (x"c3",x"48",x"d4",x"ff"),
  2454 => (x"d0",x"ff",x"78",x"ff"),
  2455 => (x"78",x"e1",x"c0",x"48"),
  2456 => (x"c1",x"48",x"d4",x"ff"),
  2457 => (x"c4",x"48",x"71",x"78"),
  2458 => (x"08",x"d4",x"ff",x"30"),
  2459 => (x"48",x"d0",x"ff",x"78"),
  2460 => (x"26",x"78",x"e0",x"c0"),
  2461 => (x"e6",x"c2",x"1e",x"4f"),
  2462 => (x"c1",x"49",x"bf",x"dc"),
  2463 => (x"c4",x"87",x"fc",x"d4"),
  2464 => (x"e8",x"48",x"d0",x"d2"),
  2465 => (x"d2",x"c4",x"78",x"bf"),
  2466 => (x"bf",x"ec",x"48",x"cc"),
  2467 => (x"d0",x"d2",x"c4",x"78"),
  2468 => (x"c3",x"49",x"4a",x"bf"),
  2469 => (x"b7",x"c8",x"99",x"ff"),
  2470 => (x"71",x"48",x"72",x"2a"),
  2471 => (x"d8",x"d2",x"c4",x"b0"),
  2472 => (x"0e",x"4f",x"26",x"58"),
  2473 => (x"5d",x"5c",x"5b",x"5e"),
  2474 => (x"ff",x"4b",x"71",x"0e"),
  2475 => (x"d2",x"c4",x"87",x"c7"),
  2476 => (x"50",x"c0",x"48",x"c8"),
  2477 => (x"de",x"e6",x"49",x"73"),
  2478 => (x"4c",x"49",x"70",x"87"),
  2479 => (x"ee",x"cb",x"9c",x"c2"),
  2480 => (x"87",x"e0",x"cb",x"49"),
  2481 => (x"d2",x"c4",x"4d",x"70"),
  2482 => (x"05",x"bf",x"97",x"c8"),
  2483 => (x"d0",x"87",x"e2",x"c1"),
  2484 => (x"d2",x"c4",x"49",x"66"),
  2485 => (x"05",x"99",x"bf",x"d4"),
  2486 => (x"66",x"d4",x"87",x"d6"),
  2487 => (x"cc",x"d2",x"c4",x"49"),
  2488 => (x"cb",x"05",x"99",x"bf"),
  2489 => (x"e5",x"49",x"73",x"87"),
  2490 => (x"98",x"70",x"87",x"ed"),
  2491 => (x"87",x"c1",x"c1",x"02"),
  2492 => (x"c0",x"fe",x"4c",x"c1"),
  2493 => (x"ca",x"49",x"75",x"87"),
  2494 => (x"98",x"70",x"87",x"f6"),
  2495 => (x"c4",x"87",x"c6",x"02"),
  2496 => (x"c1",x"48",x"c8",x"d2"),
  2497 => (x"c8",x"d2",x"c4",x"50"),
  2498 => (x"c0",x"05",x"bf",x"97"),
  2499 => (x"d2",x"c4",x"87",x"e3"),
  2500 => (x"d0",x"49",x"bf",x"d4"),
  2501 => (x"ff",x"05",x"99",x"66"),
  2502 => (x"d2",x"c4",x"87",x"d6"),
  2503 => (x"d4",x"49",x"bf",x"cc"),
  2504 => (x"ff",x"05",x"99",x"66"),
  2505 => (x"49",x"73",x"87",x"ca"),
  2506 => (x"70",x"87",x"ec",x"e4"),
  2507 => (x"ff",x"fe",x"05",x"98"),
  2508 => (x"26",x"48",x"74",x"87"),
  2509 => (x"26",x"4c",x"26",x"4d"),
  2510 => (x"0e",x"4f",x"26",x"4b"),
  2511 => (x"5d",x"5c",x"5b",x"5e"),
  2512 => (x"c0",x"86",x"f8",x"0e"),
  2513 => (x"bf",x"ec",x"4c",x"4d"),
  2514 => (x"48",x"a6",x"c4",x"7e"),
  2515 => (x"bf",x"d8",x"d2",x"c4"),
  2516 => (x"c0",x"1e",x"c1",x"78"),
  2517 => (x"fd",x"49",x"c7",x"1e"),
  2518 => (x"86",x"c8",x"87",x"c9"),
  2519 => (x"cd",x"02",x"98",x"70"),
  2520 => (x"fa",x"49",x"ff",x"87"),
  2521 => (x"da",x"c1",x"87",x"db"),
  2522 => (x"87",x"eb",x"e3",x"49"),
  2523 => (x"d2",x"c4",x"4d",x"c1"),
  2524 => (x"02",x"bf",x"97",x"c8"),
  2525 => (x"e6",x"c2",x"87",x"cf"),
  2526 => (x"c1",x"49",x"bf",x"d4"),
  2527 => (x"d8",x"e6",x"c2",x"b9"),
  2528 => (x"ce",x"fb",x"71",x"59"),
  2529 => (x"d0",x"d2",x"c4",x"87"),
  2530 => (x"e6",x"c2",x"4b",x"bf"),
  2531 => (x"c0",x"05",x"bf",x"dc"),
  2532 => (x"fd",x"c3",x"87",x"e9"),
  2533 => (x"87",x"ff",x"e2",x"49"),
  2534 => (x"e2",x"49",x"fa",x"c3"),
  2535 => (x"49",x"73",x"87",x"f9"),
  2536 => (x"71",x"99",x"ff",x"c3"),
  2537 => (x"fa",x"49",x"c0",x"1e"),
  2538 => (x"49",x"73",x"87",x"da"),
  2539 => (x"71",x"29",x"b7",x"c8"),
  2540 => (x"fa",x"49",x"c1",x"1e"),
  2541 => (x"86",x"c8",x"87",x"ce"),
  2542 => (x"c4",x"87",x"f4",x"c5"),
  2543 => (x"4b",x"bf",x"d4",x"d2"),
  2544 => (x"87",x"dd",x"02",x"9b"),
  2545 => (x"bf",x"d8",x"e6",x"c2"),
  2546 => (x"87",x"e4",x"c7",x"49"),
  2547 => (x"c4",x"05",x"98",x"70"),
  2548 => (x"d2",x"4b",x"c0",x"87"),
  2549 => (x"49",x"e0",x"c2",x"87"),
  2550 => (x"c2",x"87",x"c9",x"c7"),
  2551 => (x"c6",x"58",x"dc",x"e6"),
  2552 => (x"d8",x"e6",x"c2",x"87"),
  2553 => (x"73",x"78",x"c0",x"48"),
  2554 => (x"05",x"99",x"c2",x"49"),
  2555 => (x"eb",x"c3",x"87",x"cd"),
  2556 => (x"87",x"e3",x"e1",x"49"),
  2557 => (x"99",x"c2",x"49",x"70"),
  2558 => (x"fb",x"87",x"c2",x"02"),
  2559 => (x"c1",x"49",x"73",x"4c"),
  2560 => (x"87",x"cd",x"05",x"99"),
  2561 => (x"e1",x"49",x"f4",x"c3"),
  2562 => (x"49",x"70",x"87",x"cd"),
  2563 => (x"c2",x"02",x"99",x"c2"),
  2564 => (x"73",x"4c",x"fa",x"87"),
  2565 => (x"05",x"99",x"c8",x"49"),
  2566 => (x"f5",x"c3",x"87",x"cd"),
  2567 => (x"87",x"f7",x"e0",x"49"),
  2568 => (x"99",x"c2",x"49",x"70"),
  2569 => (x"c4",x"87",x"d5",x"02"),
  2570 => (x"02",x"bf",x"dc",x"d2"),
  2571 => (x"c1",x"48",x"87",x"ca"),
  2572 => (x"e0",x"d2",x"c4",x"88"),
  2573 => (x"87",x"c2",x"c0",x"58"),
  2574 => (x"4d",x"c1",x"4c",x"ff"),
  2575 => (x"99",x"c4",x"49",x"73"),
  2576 => (x"c3",x"87",x"cd",x"05"),
  2577 => (x"ce",x"e0",x"49",x"f2"),
  2578 => (x"c2",x"49",x"70",x"87"),
  2579 => (x"87",x"dc",x"02",x"99"),
  2580 => (x"bf",x"dc",x"d2",x"c4"),
  2581 => (x"b7",x"c7",x"48",x"7e"),
  2582 => (x"cb",x"c0",x"03",x"a8"),
  2583 => (x"c1",x"48",x"6e",x"87"),
  2584 => (x"e0",x"d2",x"c4",x"80"),
  2585 => (x"87",x"c2",x"c0",x"58"),
  2586 => (x"4d",x"c1",x"4c",x"fe"),
  2587 => (x"ff",x"49",x"fd",x"c3"),
  2588 => (x"70",x"87",x"e4",x"df"),
  2589 => (x"02",x"99",x"c2",x"49"),
  2590 => (x"d2",x"c4",x"87",x"d5"),
  2591 => (x"c0",x"02",x"bf",x"dc"),
  2592 => (x"d2",x"c4",x"87",x"c9"),
  2593 => (x"78",x"c0",x"48",x"dc"),
  2594 => (x"fd",x"87",x"c2",x"c0"),
  2595 => (x"c3",x"4d",x"c1",x"4c"),
  2596 => (x"df",x"ff",x"49",x"fa"),
  2597 => (x"49",x"70",x"87",x"c1"),
  2598 => (x"c0",x"02",x"99",x"c2"),
  2599 => (x"d2",x"c4",x"87",x"d9"),
  2600 => (x"c7",x"48",x"bf",x"dc"),
  2601 => (x"c0",x"03",x"a8",x"b7"),
  2602 => (x"d2",x"c4",x"87",x"c9"),
  2603 => (x"78",x"c7",x"48",x"dc"),
  2604 => (x"fc",x"87",x"c2",x"c0"),
  2605 => (x"c0",x"4d",x"c1",x"4c"),
  2606 => (x"c0",x"03",x"ac",x"b7"),
  2607 => (x"66",x"c4",x"87",x"d3"),
  2608 => (x"80",x"e0",x"c1",x"48"),
  2609 => (x"bf",x"6e",x"7e",x"70"),
  2610 => (x"87",x"c5",x"c0",x"02"),
  2611 => (x"73",x"49",x"74",x"4b"),
  2612 => (x"c3",x"1e",x"c0",x"0f"),
  2613 => (x"da",x"c1",x"1e",x"f0"),
  2614 => (x"87",x"c7",x"f7",x"49"),
  2615 => (x"98",x"70",x"86",x"c8"),
  2616 => (x"87",x"d8",x"c0",x"02"),
  2617 => (x"bf",x"dc",x"d2",x"c4"),
  2618 => (x"cc",x"49",x"6e",x"7e"),
  2619 => (x"4a",x"66",x"c4",x"91"),
  2620 => (x"02",x"6a",x"82",x"71"),
  2621 => (x"4b",x"87",x"c5",x"c0"),
  2622 => (x"0f",x"73",x"49",x"6e"),
  2623 => (x"c0",x"02",x"9d",x"75"),
  2624 => (x"d2",x"c4",x"87",x"c8"),
  2625 => (x"f2",x"49",x"bf",x"dc"),
  2626 => (x"e6",x"c2",x"87",x"d6"),
  2627 => (x"c0",x"02",x"bf",x"e0"),
  2628 => (x"c2",x"49",x"87",x"dd"),
  2629 => (x"98",x"70",x"87",x"da"),
  2630 => (x"87",x"d3",x"c0",x"02"),
  2631 => (x"bf",x"dc",x"d2",x"c4"),
  2632 => (x"87",x"fc",x"f1",x"49"),
  2633 => (x"d8",x"f3",x"49",x"c0"),
  2634 => (x"e0",x"e6",x"c2",x"87"),
  2635 => (x"f8",x"78",x"c0",x"48"),
  2636 => (x"26",x"4d",x"26",x"8e"),
  2637 => (x"26",x"4b",x"26",x"4c"),
  2638 => (x"5b",x"5e",x"0e",x"4f"),
  2639 => (x"fc",x"0e",x"5d",x"5c"),
  2640 => (x"c4",x"4c",x"71",x"86"),
  2641 => (x"49",x"bf",x"d8",x"d2"),
  2642 => (x"4d",x"a1",x"d4",x"c1"),
  2643 => (x"69",x"81",x"d8",x"c1"),
  2644 => (x"02",x"9c",x"74",x"7e"),
  2645 => (x"a5",x"c4",x"87",x"cf"),
  2646 => (x"c4",x"7b",x"74",x"4b"),
  2647 => (x"49",x"bf",x"d8",x"d2"),
  2648 => (x"6e",x"87",x"cb",x"f2"),
  2649 => (x"05",x"9c",x"74",x"7b"),
  2650 => (x"4b",x"c0",x"87",x"c4"),
  2651 => (x"4b",x"c1",x"87",x"c2"),
  2652 => (x"cc",x"f2",x"49",x"73"),
  2653 => (x"02",x"66",x"d4",x"87"),
  2654 => (x"c0",x"49",x"87",x"c8"),
  2655 => (x"4a",x"70",x"87",x"e6"),
  2656 => (x"4a",x"c0",x"87",x"c2"),
  2657 => (x"5a",x"e4",x"e6",x"c2"),
  2658 => (x"4d",x"26",x"8e",x"fc"),
  2659 => (x"4b",x"26",x"4c",x"26"),
  2660 => (x"00",x"00",x"4f",x"26"),
  2661 => (x"00",x"00",x"00",x"00"),
  2662 => (x"00",x"00",x"00",x"00"),
  2663 => (x"00",x"00",x"00",x"00"),
  2664 => (x"00",x"00",x"00",x"00"),
  2665 => (x"ff",x"4a",x"71",x"1e"),
  2666 => (x"72",x"49",x"bf",x"c8"),
  2667 => (x"4f",x"26",x"48",x"a1"),
  2668 => (x"bf",x"c8",x"ff",x"1e"),
  2669 => (x"c0",x"c0",x"fe",x"89"),
  2670 => (x"a9",x"c0",x"c0",x"c0"),
  2671 => (x"c0",x"87",x"c4",x"01"),
  2672 => (x"c1",x"87",x"c2",x"4a"),
  2673 => (x"26",x"48",x"72",x"4a"),
  2674 => (x"5b",x"5e",x"0e",x"4f"),
  2675 => (x"71",x"0e",x"5d",x"5c"),
  2676 => (x"4c",x"d4",x"ff",x"4b"),
  2677 => (x"c0",x"48",x"66",x"d0"),
  2678 => (x"ff",x"49",x"d6",x"78"),
  2679 => (x"c3",x"87",x"f5",x"db"),
  2680 => (x"49",x"6c",x"7c",x"ff"),
  2681 => (x"71",x"99",x"ff",x"c3"),
  2682 => (x"f0",x"c3",x"49",x"4d"),
  2683 => (x"a9",x"e0",x"c1",x"99"),
  2684 => (x"c3",x"87",x"cb",x"05"),
  2685 => (x"48",x"6c",x"7c",x"ff"),
  2686 => (x"66",x"d0",x"98",x"c3"),
  2687 => (x"ff",x"c3",x"78",x"08"),
  2688 => (x"49",x"4a",x"6c",x"7c"),
  2689 => (x"ff",x"c3",x"31",x"c8"),
  2690 => (x"71",x"4a",x"6c",x"7c"),
  2691 => (x"c8",x"49",x"72",x"b2"),
  2692 => (x"7c",x"ff",x"c3",x"31"),
  2693 => (x"b2",x"71",x"4a",x"6c"),
  2694 => (x"31",x"c8",x"49",x"72"),
  2695 => (x"6c",x"7c",x"ff",x"c3"),
  2696 => (x"ff",x"b2",x"71",x"4a"),
  2697 => (x"e0",x"c0",x"48",x"d0"),
  2698 => (x"02",x"9b",x"73",x"78"),
  2699 => (x"7b",x"72",x"87",x"c2"),
  2700 => (x"4d",x"26",x"48",x"75"),
  2701 => (x"4b",x"26",x"4c",x"26"),
  2702 => (x"26",x"1e",x"4f",x"26"),
  2703 => (x"5b",x"5e",x"0e",x"4f"),
  2704 => (x"86",x"f8",x"0e",x"5c"),
  2705 => (x"a6",x"c8",x"1e",x"76"),
  2706 => (x"87",x"fd",x"fd",x"49"),
  2707 => (x"4b",x"70",x"86",x"c4"),
  2708 => (x"a8",x"c4",x"48",x"6e"),
  2709 => (x"87",x"f4",x"c2",x"03"),
  2710 => (x"f0",x"c3",x"4a",x"73"),
  2711 => (x"aa",x"d0",x"c1",x"9a"),
  2712 => (x"c1",x"87",x"c7",x"02"),
  2713 => (x"c2",x"05",x"aa",x"e0"),
  2714 => (x"49",x"73",x"87",x"e2"),
  2715 => (x"c3",x"02",x"99",x"c8"),
  2716 => (x"87",x"c6",x"ff",x"87"),
  2717 => (x"9c",x"c3",x"4c",x"73"),
  2718 => (x"c1",x"05",x"ac",x"c2"),
  2719 => (x"66",x"c4",x"87",x"c4"),
  2720 => (x"71",x"31",x"c9",x"49"),
  2721 => (x"4a",x"66",x"c4",x"1e"),
  2722 => (x"c4",x"92",x"c8",x"c1"),
  2723 => (x"72",x"49",x"e0",x"d2"),
  2724 => (x"f7",x"c3",x"fe",x"81"),
  2725 => (x"ff",x"49",x"d8",x"87"),
  2726 => (x"c8",x"87",x"f9",x"d8"),
  2727 => (x"ff",x"c3",x"1e",x"c0"),
  2728 => (x"db",x"fd",x"49",x"e0"),
  2729 => (x"d0",x"ff",x"87",x"c1"),
  2730 => (x"78",x"e0",x"c0",x"48"),
  2731 => (x"1e",x"e0",x"ff",x"c3"),
  2732 => (x"c1",x"4a",x"66",x"cc"),
  2733 => (x"d2",x"c4",x"92",x"c8"),
  2734 => (x"81",x"72",x"49",x"e0"),
  2735 => (x"87",x"c6",x"ff",x"fd"),
  2736 => (x"ac",x"c1",x"86",x"cc"),
  2737 => (x"87",x"c4",x"c1",x"05"),
  2738 => (x"c9",x"49",x"66",x"c4"),
  2739 => (x"c4",x"1e",x"71",x"31"),
  2740 => (x"c8",x"c1",x"4a",x"66"),
  2741 => (x"e0",x"d2",x"c4",x"92"),
  2742 => (x"fe",x"81",x"72",x"49"),
  2743 => (x"c3",x"87",x"ed",x"c2"),
  2744 => (x"c8",x"1e",x"e0",x"ff"),
  2745 => (x"c8",x"c1",x"4a",x"66"),
  2746 => (x"e0",x"d2",x"c4",x"92"),
  2747 => (x"fd",x"81",x"72",x"49"),
  2748 => (x"d7",x"87",x"c4",x"fd"),
  2749 => (x"db",x"d7",x"ff",x"49"),
  2750 => (x"1e",x"c0",x"c8",x"87"),
  2751 => (x"49",x"e0",x"ff",x"c3"),
  2752 => (x"87",x"c0",x"d9",x"fd"),
  2753 => (x"d0",x"ff",x"86",x"cc"),
  2754 => (x"78",x"e0",x"c0",x"48"),
  2755 => (x"4c",x"26",x"8e",x"f8"),
  2756 => (x"4f",x"26",x"4b",x"26"),
  2757 => (x"5c",x"5b",x"5e",x"0e"),
  2758 => (x"4a",x"71",x"0e",x"5d"),
  2759 => (x"d0",x"4c",x"d4",x"ff"),
  2760 => (x"b7",x"c3",x"4d",x"66"),
  2761 => (x"87",x"c5",x"06",x"ad"),
  2762 => (x"e2",x"c1",x"48",x"c0"),
  2763 => (x"75",x"1e",x"72",x"87"),
  2764 => (x"93",x"c8",x"c1",x"4b"),
  2765 => (x"83",x"e0",x"d2",x"c4"),
  2766 => (x"f5",x"fd",x"49",x"73"),
  2767 => (x"83",x"c8",x"87",x"f5"),
  2768 => (x"d0",x"ff",x"4b",x"6b"),
  2769 => (x"78",x"e1",x"c8",x"48"),
  2770 => (x"48",x"73",x"7c",x"dd"),
  2771 => (x"70",x"98",x"ff",x"c3"),
  2772 => (x"c8",x"49",x"73",x"7c"),
  2773 => (x"48",x"71",x"29",x"b7"),
  2774 => (x"70",x"98",x"ff",x"c3"),
  2775 => (x"d0",x"49",x"73",x"7c"),
  2776 => (x"48",x"71",x"29",x"b7"),
  2777 => (x"70",x"98",x"ff",x"c3"),
  2778 => (x"d8",x"48",x"73",x"7c"),
  2779 => (x"7c",x"70",x"28",x"b7"),
  2780 => (x"7c",x"7c",x"7c",x"c0"),
  2781 => (x"7c",x"7c",x"7c",x"7c"),
  2782 => (x"7c",x"7c",x"7c",x"7c"),
  2783 => (x"48",x"d0",x"ff",x"7c"),
  2784 => (x"75",x"78",x"e0",x"c0"),
  2785 => (x"ff",x"49",x"dc",x"1e"),
  2786 => (x"c8",x"87",x"ee",x"d5"),
  2787 => (x"26",x"48",x"73",x"86"),
  2788 => (x"26",x"4c",x"26",x"4d"),
  2789 => (x"1e",x"4f",x"26",x"4b"),
  2790 => (x"86",x"fc",x"1e",x"73"),
  2791 => (x"f0",x"c0",x"4b",x"71"),
  2792 => (x"ec",x"c0",x"4a",x"a3"),
  2793 => (x"82",x"69",x"49",x"a3"),
  2794 => (x"69",x"52",x"66",x"cc"),
  2795 => (x"70",x"80",x"c1",x"48"),
  2796 => (x"98",x"cf",x"48",x"7e"),
  2797 => (x"8e",x"fc",x"79",x"70"),
  2798 => (x"4f",x"26",x"4b",x"26"),
  2799 => (x"5c",x"5b",x"5e",x"0e"),
  2800 => (x"e9",x"4b",x"71",x"0e"),
  2801 => (x"4c",x"70",x"87",x"f6"),
  2802 => (x"87",x"fc",x"c6",x"ff"),
  2803 => (x"c2",x"49",x"66",x"cc"),
  2804 => (x"dc",x"02",x"99",x"c0"),
  2805 => (x"05",x"9c",x"74",x"87"),
  2806 => (x"e0",x"c3",x"87",x"ca"),
  2807 => (x"fe",x"49",x"73",x"1e"),
  2808 => (x"86",x"c4",x"87",x"f5"),
  2809 => (x"c4",x"1e",x"e0",x"c3"),
  2810 => (x"ff",x"49",x"cc",x"d1"),
  2811 => (x"c4",x"87",x"ff",x"c9"),
  2812 => (x"49",x"66",x"cc",x"86"),
  2813 => (x"02",x"99",x"c0",x"c4"),
  2814 => (x"9c",x"74",x"87",x"dc"),
  2815 => (x"c3",x"87",x"ca",x"05"),
  2816 => (x"49",x"73",x"1e",x"f0"),
  2817 => (x"c4",x"87",x"d0",x"fe"),
  2818 => (x"1e",x"f0",x"c3",x"86"),
  2819 => (x"49",x"cc",x"d1",x"c4"),
  2820 => (x"87",x"da",x"c9",x"ff"),
  2821 => (x"9c",x"74",x"86",x"c4"),
  2822 => (x"cc",x"87",x"cf",x"05"),
  2823 => (x"ff",x"c1",x"49",x"66"),
  2824 => (x"73",x"1e",x"71",x"99"),
  2825 => (x"87",x"ef",x"fd",x"49"),
  2826 => (x"66",x"cc",x"86",x"c4"),
  2827 => (x"99",x"ff",x"c1",x"49"),
  2828 => (x"d1",x"c4",x"1e",x"71"),
  2829 => (x"c8",x"ff",x"49",x"cc"),
  2830 => (x"c5",x"ff",x"87",x"f4"),
  2831 => (x"8e",x"fc",x"87",x"c2"),
  2832 => (x"4b",x"26",x"4c",x"26"),
  2833 => (x"5e",x"0e",x"4f",x"26"),
  2834 => (x"fc",x"0e",x"5c",x"5b"),
  2835 => (x"f7",x"c4",x"ff",x"86"),
  2836 => (x"c8",x"f3",x"c2",x"87"),
  2837 => (x"d7",x"f5",x"49",x"bf"),
  2838 => (x"02",x"98",x"70",x"87"),
  2839 => (x"c4",x"87",x"dc",x"c1"),
  2840 => (x"48",x"bf",x"ec",x"d7"),
  2841 => (x"bf",x"f0",x"d7",x"c4"),
  2842 => (x"ce",x"c1",x"02",x"a8"),
  2843 => (x"f4",x"d7",x"c4",x"87"),
  2844 => (x"ec",x"d7",x"c4",x"49"),
  2845 => (x"4c",x"11",x"81",x"bf"),
  2846 => (x"aa",x"e0",x"c3",x"4a"),
  2847 => (x"c3",x"87",x"c6",x"02"),
  2848 => (x"c4",x"05",x"aa",x"f0"),
  2849 => (x"c2",x"4b",x"c4",x"87"),
  2850 => (x"73",x"4b",x"cf",x"87"),
  2851 => (x"87",x"d4",x"f4",x"49"),
  2852 => (x"58",x"cc",x"f3",x"c2"),
  2853 => (x"c8",x"48",x"d0",x"ff"),
  2854 => (x"d4",x"ff",x"78",x"e1"),
  2855 => (x"74",x"78",x"c5",x"48"),
  2856 => (x"08",x"d4",x"ff",x"48"),
  2857 => (x"48",x"d0",x"ff",x"78"),
  2858 => (x"c4",x"78",x"e0",x"c0"),
  2859 => (x"48",x"bf",x"ec",x"d7"),
  2860 => (x"7e",x"70",x"80",x"c1"),
  2861 => (x"c4",x"98",x"cf",x"48"),
  2862 => (x"ff",x"58",x"f0",x"d7"),
  2863 => (x"fc",x"87",x"c1",x"c3"),
  2864 => (x"26",x"4c",x"26",x"8e"),
  2865 => (x"00",x"4f",x"26",x"4b"),
  2866 => (x"00",x"00",x"00",x"00"),
  2867 => (x"5c",x"5b",x"5e",x"0e"),
  2868 => (x"dc",x"ff",x"0e",x"5d"),
  2869 => (x"c4",x"7e",x"c0",x"86"),
  2870 => (x"49",x"bf",x"c8",x"d7"),
  2871 => (x"1e",x"71",x"81",x"c2"),
  2872 => (x"4a",x"c6",x"1e",x"72"),
  2873 => (x"87",x"eb",x"d0",x"fd"),
  2874 => (x"4a",x"26",x"48",x"71"),
  2875 => (x"a6",x"cc",x"49",x"26"),
  2876 => (x"c8",x"d7",x"c4",x"58"),
  2877 => (x"81",x"c4",x"49",x"bf"),
  2878 => (x"1e",x"72",x"1e",x"71"),
  2879 => (x"d0",x"fd",x"4a",x"c6"),
  2880 => (x"48",x"71",x"87",x"d1"),
  2881 => (x"49",x"26",x"4a",x"26"),
  2882 => (x"fc",x"58",x"a6",x"d0"),
  2883 => (x"fe",x"c2",x"87",x"f8"),
  2884 => (x"f2",x"49",x"bf",x"dc"),
  2885 => (x"98",x"70",x"87",x"da"),
  2886 => (x"87",x"f2",x"c9",x"02"),
  2887 => (x"f2",x"49",x"e0",x"c0"),
  2888 => (x"fe",x"c2",x"87",x"c2"),
  2889 => (x"4c",x"c0",x"58",x"e0"),
  2890 => (x"91",x"c4",x"49",x"74"),
  2891 => (x"69",x"81",x"d0",x"fe"),
  2892 => (x"c4",x"49",x"74",x"4a"),
  2893 => (x"81",x"bf",x"c8",x"d7"),
  2894 => (x"d7",x"c4",x"91",x"c4"),
  2895 => (x"79",x"72",x"81",x"d4"),
  2896 => (x"87",x"d2",x"02",x"9a"),
  2897 => (x"89",x"c1",x"49",x"72"),
  2898 => (x"48",x"6e",x"9a",x"71"),
  2899 => (x"7e",x"70",x"80",x"c1"),
  2900 => (x"ff",x"05",x"9a",x"72"),
  2901 => (x"84",x"c1",x"87",x"ee"),
  2902 => (x"04",x"ac",x"b7",x"c2"),
  2903 => (x"6e",x"87",x"c9",x"ff"),
  2904 => (x"b7",x"fc",x"c0",x"48"),
  2905 => (x"e5",x"c8",x"04",x"a8"),
  2906 => (x"74",x"4c",x"c0",x"87"),
  2907 => (x"82",x"66",x"c8",x"4a"),
  2908 => (x"d7",x"c4",x"92",x"c4"),
  2909 => (x"49",x"74",x"82",x"d4"),
  2910 => (x"c4",x"81",x"66",x"cc"),
  2911 => (x"d4",x"d7",x"c4",x"91"),
  2912 => (x"69",x"4a",x"6a",x"81"),
  2913 => (x"74",x"b9",x"72",x"49"),
  2914 => (x"c8",x"d7",x"c4",x"4b"),
  2915 => (x"93",x"c4",x"83",x"bf"),
  2916 => (x"83",x"d4",x"d7",x"c4"),
  2917 => (x"48",x"72",x"ba",x"6b"),
  2918 => (x"a6",x"d8",x"98",x"71"),
  2919 => (x"c4",x"49",x"74",x"58"),
  2920 => (x"81",x"bf",x"c8",x"d7"),
  2921 => (x"d7",x"c4",x"91",x"c4"),
  2922 => (x"7e",x"69",x"81",x"d4"),
  2923 => (x"c0",x"48",x"a6",x"d8"),
  2924 => (x"5c",x"a6",x"d4",x"78"),
  2925 => (x"df",x"49",x"66",x"d4"),
  2926 => (x"e0",x"c6",x"02",x"29"),
  2927 => (x"4a",x"66",x"d0",x"87"),
  2928 => (x"d8",x"92",x"e0",x"c0"),
  2929 => (x"ff",x"c0",x"82",x"66"),
  2930 => (x"70",x"88",x"72",x"48"),
  2931 => (x"48",x"a6",x"dc",x"4a"),
  2932 => (x"80",x"c4",x"78",x"c0"),
  2933 => (x"4c",x"6e",x"78",x"c0"),
  2934 => (x"d7",x"c4",x"2c",x"df"),
  2935 => (x"78",x"c1",x"48",x"c4"),
  2936 => (x"31",x"c3",x"49",x"72"),
  2937 => (x"b1",x"72",x"2a",x"b7"),
  2938 => (x"c4",x"99",x"ff",x"c0"),
  2939 => (x"d8",x"f0",x"c3",x"91"),
  2940 => (x"6d",x"85",x"71",x"4d"),
  2941 => (x"c0",x"c4",x"49",x"4b"),
  2942 => (x"d6",x"02",x"99",x"c0"),
  2943 => (x"02",x"9c",x"74",x"87"),
  2944 => (x"c8",x"87",x"c7",x"c0"),
  2945 => (x"c5",x"78",x"c0",x"80"),
  2946 => (x"d7",x"c4",x"87",x"d3"),
  2947 => (x"78",x"c1",x"48",x"cc"),
  2948 => (x"74",x"87",x"ca",x"c5"),
  2949 => (x"87",x"d8",x"02",x"9c"),
  2950 => (x"c0",x"c2",x"49",x"73"),
  2951 => (x"c0",x"02",x"99",x"c0"),
  2952 => (x"b7",x"d0",x"87",x"c3"),
  2953 => (x"fd",x"48",x"6d",x"2b"),
  2954 => (x"70",x"98",x"ff",x"ff"),
  2955 => (x"87",x"f8",x"c0",x"7d"),
  2956 => (x"bf",x"cc",x"d7",x"c4"),
  2957 => (x"87",x"f0",x"c0",x"02"),
  2958 => (x"b7",x"d0",x"48",x"73"),
  2959 => (x"58",x"a6",x"c8",x"28"),
  2960 => (x"c0",x"02",x"98",x"70"),
  2961 => (x"d7",x"c4",x"87",x"e2"),
  2962 => (x"c0",x"49",x"bf",x"d0"),
  2963 => (x"02",x"99",x"c0",x"e0"),
  2964 => (x"70",x"87",x"ca",x"c0"),
  2965 => (x"c0",x"e0",x"c0",x"49"),
  2966 => (x"cb",x"c0",x"02",x"99"),
  2967 => (x"c2",x"48",x"6d",x"87"),
  2968 => (x"70",x"b0",x"c0",x"c0"),
  2969 => (x"4b",x"66",x"c4",x"7d"),
  2970 => (x"c0",x"c8",x"49",x"73"),
  2971 => (x"c2",x"02",x"99",x"c0"),
  2972 => (x"d7",x"c4",x"87",x"c9"),
  2973 => (x"cc",x"4a",x"bf",x"d0"),
  2974 => (x"c0",x"02",x"9a",x"c0"),
  2975 => (x"c0",x"c4",x"87",x"cf"),
  2976 => (x"d8",x"c0",x"02",x"8a"),
  2977 => (x"c0",x"02",x"8a",x"87"),
  2978 => (x"df",x"c1",x"87",x"fa"),
  2979 => (x"c3",x"49",x"73",x"87"),
  2980 => (x"91",x"c2",x"99",x"ff"),
  2981 => (x"81",x"cc",x"f0",x"c3"),
  2982 => (x"de",x"c1",x"4b",x"11"),
  2983 => (x"c3",x"49",x"73",x"87"),
  2984 => (x"91",x"c2",x"99",x"ff"),
  2985 => (x"81",x"cc",x"f0",x"c3"),
  2986 => (x"4b",x"11",x"81",x"c1"),
  2987 => (x"c0",x"02",x"9c",x"74"),
  2988 => (x"e0",x"c0",x"87",x"c9"),
  2989 => (x"78",x"d2",x"48",x"a6"),
  2990 => (x"dc",x"87",x"c0",x"c1"),
  2991 => (x"d2",x"c4",x"48",x"a6"),
  2992 => (x"87",x"f7",x"c0",x"78"),
  2993 => (x"ff",x"c3",x"49",x"73"),
  2994 => (x"c3",x"91",x"c2",x"99"),
  2995 => (x"c1",x"81",x"cc",x"f0"),
  2996 => (x"74",x"4b",x"11",x"81"),
  2997 => (x"ca",x"c0",x"02",x"9c"),
  2998 => (x"a6",x"e0",x"c0",x"87"),
  2999 => (x"78",x"d9",x"c1",x"48"),
  3000 => (x"dc",x"87",x"d8",x"c0"),
  3001 => (x"d9",x"c5",x"48",x"a6"),
  3002 => (x"87",x"cf",x"c0",x"78"),
  3003 => (x"ff",x"c3",x"49",x"73"),
  3004 => (x"c3",x"91",x"c2",x"99"),
  3005 => (x"c1",x"81",x"cc",x"f0"),
  3006 => (x"74",x"4b",x"11",x"81"),
  3007 => (x"dc",x"c0",x"02",x"9c"),
  3008 => (x"ff",x"49",x"73",x"87"),
  3009 => (x"c0",x"fc",x"c7",x"b9"),
  3010 => (x"c4",x"48",x"71",x"99"),
  3011 => (x"98",x"bf",x"d0",x"d7"),
  3012 => (x"58",x"d4",x"d7",x"c4"),
  3013 => (x"c4",x"9b",x"ff",x"c3"),
  3014 => (x"d4",x"c0",x"b3",x"c0"),
  3015 => (x"c7",x"49",x"73",x"87"),
  3016 => (x"71",x"99",x"c0",x"fc"),
  3017 => (x"d0",x"d7",x"c4",x"48"),
  3018 => (x"d7",x"c4",x"b0",x"bf"),
  3019 => (x"ff",x"c3",x"58",x"d4"),
  3020 => (x"02",x"66",x"dc",x"9b"),
  3021 => (x"1e",x"87",x"ca",x"c0"),
  3022 => (x"49",x"c4",x"d7",x"c4"),
  3023 => (x"c4",x"87",x"fd",x"f1"),
  3024 => (x"c4",x"1e",x"73",x"86"),
  3025 => (x"f1",x"49",x"c4",x"d7"),
  3026 => (x"86",x"c4",x"87",x"f2"),
  3027 => (x"02",x"66",x"e0",x"c0"),
  3028 => (x"1e",x"87",x"ca",x"c0"),
  3029 => (x"49",x"c4",x"d7",x"c4"),
  3030 => (x"c4",x"87",x"e1",x"f1"),
  3031 => (x"48",x"66",x"d4",x"86"),
  3032 => (x"a6",x"d8",x"30",x"c1"),
  3033 => (x"c1",x"48",x"6e",x"58"),
  3034 => (x"d8",x"7e",x"70",x"30"),
  3035 => (x"80",x"c1",x"48",x"66"),
  3036 => (x"c0",x"58",x"a6",x"dc"),
  3037 => (x"04",x"a8",x"b7",x"e0"),
  3038 => (x"d0",x"87",x"f9",x"f8"),
  3039 => (x"84",x"c1",x"4c",x"66"),
  3040 => (x"04",x"ac",x"b7",x"c2"),
  3041 => (x"c4",x"87",x"e4",x"f7"),
  3042 => (x"c8",x"48",x"c8",x"d7"),
  3043 => (x"dc",x"ff",x"78",x"66"),
  3044 => (x"26",x"4d",x"26",x"8e"),
  3045 => (x"26",x"4b",x"26",x"4c"),
  3046 => (x"00",x"00",x"00",x"4f"),
  3047 => (x"00",x"00",x"00",x"00"),
  3048 => (x"72",x"4a",x"c0",x"1e"),
  3049 => (x"c4",x"91",x"c4",x"49"),
  3050 => (x"ff",x"81",x"d4",x"d7"),
  3051 => (x"c6",x"82",x"c1",x"79"),
  3052 => (x"ee",x"04",x"aa",x"b7"),
  3053 => (x"c8",x"d7",x"c4",x"87"),
  3054 => (x"40",x"40",x"c0",x"48"),
  3055 => (x"0e",x"4f",x"26",x"78"),
  3056 => (x"0e",x"5c",x"5b",x"5e"),
  3057 => (x"d4",x"ff",x"4a",x"71"),
  3058 => (x"4b",x"66",x"cc",x"4c"),
  3059 => (x"c8",x"48",x"d0",x"ff"),
  3060 => (x"7c",x"c2",x"78",x"c5"),
  3061 => (x"8b",x"c1",x"49",x"73"),
  3062 => (x"cd",x"02",x"99",x"71"),
  3063 => (x"12",x"7c",x"12",x"87"),
  3064 => (x"c1",x"49",x"73",x"7c"),
  3065 => (x"05",x"99",x"71",x"8b"),
  3066 => (x"d0",x"ff",x"87",x"f3"),
  3067 => (x"26",x"78",x"c4",x"48"),
  3068 => (x"26",x"4b",x"26",x"4c"),
  3069 => (x"4a",x"71",x"1e",x"4f"),
  3070 => (x"c8",x"48",x"d0",x"ff"),
  3071 => (x"d4",x"ff",x"78",x"c5"),
  3072 => (x"c8",x"78",x"c3",x"48"),
  3073 => (x"49",x"72",x"1e",x"c0"),
  3074 => (x"87",x"db",x"c5",x"fd"),
  3075 => (x"c4",x"48",x"d0",x"ff"),
  3076 => (x"26",x"8e",x"fc",x"78"),
  3077 => (x"d0",x"ff",x"1e",x"4f"),
  3078 => (x"78",x"c5",x"c8",x"48"),
  3079 => (x"c6",x"48",x"d4",x"ff"),
  3080 => (x"ff",x"48",x"71",x"78"),
  3081 => (x"ff",x"78",x"08",x"d4"),
  3082 => (x"78",x"c4",x"48",x"d0"),
  3083 => (x"ff",x"1e",x"4f",x"26"),
  3084 => (x"c5",x"c8",x"48",x"d0"),
  3085 => (x"48",x"d4",x"ff",x"78"),
  3086 => (x"d0",x"ff",x"78",x"ca"),
  3087 => (x"26",x"78",x"c4",x"48"),
  3088 => (x"5b",x"5e",x"0e",x"4f"),
  3089 => (x"ff",x"0e",x"5d",x"5c"),
  3090 => (x"7e",x"71",x"86",x"d4"),
  3091 => (x"81",x"ca",x"49",x"6e"),
  3092 => (x"48",x"49",x"69",x"97"),
  3093 => (x"d4",x"28",x"b7",x"c5"),
  3094 => (x"49",x"6e",x"58",x"a6"),
  3095 => (x"69",x"97",x"81",x"c1"),
  3096 => (x"b7",x"c5",x"48",x"49"),
  3097 => (x"58",x"a6",x"d8",x"28"),
  3098 => (x"48",x"bf",x"97",x"6e"),
  3099 => (x"df",x"58",x"a6",x"dc"),
  3100 => (x"c0",x"c0",x"d0",x"99"),
  3101 => (x"c2",x"4a",x"6e",x"91"),
  3102 => (x"c0",x"48",x"12",x"82"),
  3103 => (x"70",x"58",x"a6",x"e0"),
  3104 => (x"92",x"c0",x"c4",x"4a"),
  3105 => (x"6e",x"49",x"a1",x"72"),
  3106 => (x"12",x"82",x"c3",x"4a"),
  3107 => (x"a6",x"e4",x"c0",x"48"),
  3108 => (x"c0",x"80",x"71",x"58"),
  3109 => (x"6e",x"58",x"a6",x"e8"),
  3110 => (x"c8",x"80",x"c4",x"48"),
  3111 => (x"66",x"c4",x"58",x"a6"),
  3112 => (x"9c",x"4c",x"bf",x"97"),
  3113 => (x"c4",x"87",x"c3",x"05"),
  3114 => (x"66",x"d0",x"4c",x"c0"),
  3115 => (x"a8",x"b7",x"c2",x"48"),
  3116 => (x"87",x"f1",x"cf",x"03"),
  3117 => (x"c1",x"49",x"66",x"d0"),
  3118 => (x"d4",x"c4",x"91",x"c8"),
  3119 => (x"80",x"71",x"48",x"f0"),
  3120 => (x"cc",x"58",x"a6",x"d0"),
  3121 => (x"80",x"c8",x"48",x"66"),
  3122 => (x"c8",x"58",x"a6",x"cc"),
  3123 => (x"cf",x"02",x"bf",x"66"),
  3124 => (x"c9",x"48",x"87",x"d3"),
  3125 => (x"a6",x"ec",x"c0",x"28"),
  3126 => (x"02",x"66",x"d8",x"58"),
  3127 => (x"4d",x"87",x"e3",x"c2"),
  3128 => (x"c3",x"02",x"8d",x"c3"),
  3129 => (x"8d",x"c1",x"87",x"c3"),
  3130 => (x"87",x"d6",x"c2",x"02"),
  3131 => (x"c4",x"02",x"8d",x"c4"),
  3132 => (x"8d",x"c2",x"87",x"cf"),
  3133 => (x"87",x"d6",x"c7",x"02"),
  3134 => (x"ca",x"02",x"8d",x"c8"),
  3135 => (x"02",x"8d",x"87",x"e5"),
  3136 => (x"cb",x"87",x"e6",x"cc"),
  3137 => (x"87",x"cf",x"02",x"8d"),
  3138 => (x"c3",x"02",x"8d",x"c3"),
  3139 => (x"8d",x"c2",x"87",x"f3"),
  3140 => (x"87",x"fa",x"c6",x"02"),
  3141 => (x"d4",x"87",x"fc",x"cd"),
  3142 => (x"d3",x"c1",x"05",x"66"),
  3143 => (x"e0",x"ff",x"c3",x"87"),
  3144 => (x"c8",x"4a",x"c0",x"4b"),
  3145 => (x"fe",x"fc",x"49",x"c0"),
  3146 => (x"e8",x"c0",x"87",x"e8"),
  3147 => (x"89",x"c1",x"49",x"66"),
  3148 => (x"2a",x"d8",x"4a",x"71"),
  3149 => (x"97",x"e4",x"ff",x"c3"),
  3150 => (x"d0",x"4a",x"71",x"5a"),
  3151 => (x"e5",x"ff",x"c3",x"2a"),
  3152 => (x"4a",x"71",x"5a",x"97"),
  3153 => (x"ff",x"c3",x"2a",x"c8"),
  3154 => (x"c3",x"5a",x"97",x"e6"),
  3155 => (x"59",x"97",x"e7",x"ff"),
  3156 => (x"c2",x"80",x"c3",x"48"),
  3157 => (x"f9",x"1e",x"c4",x"50"),
  3158 => (x"e2",x"f9",x"49",x"a0"),
  3159 => (x"c0",x"86",x"c4",x"87"),
  3160 => (x"87",x"f1",x"fa",x"49"),
  3161 => (x"49",x"e8",x"d3",x"c3"),
  3162 => (x"c0",x"81",x"66",x"d0"),
  3163 => (x"87",x"f8",x"cc",x"51"),
  3164 => (x"e0",x"fa",x"49",x"c2"),
  3165 => (x"e8",x"d3",x"c3",x"87"),
  3166 => (x"81",x"66",x"d0",x"49"),
  3167 => (x"cc",x"51",x"e5",x"c0"),
  3168 => (x"66",x"d4",x"87",x"e6"),
  3169 => (x"c3",x"87",x"d0",x"05"),
  3170 => (x"d0",x"49",x"e8",x"d3"),
  3171 => (x"51",x"c0",x"81",x"66"),
  3172 => (x"87",x"c1",x"fa",x"49"),
  3173 => (x"c3",x"87",x"d1",x"cc"),
  3174 => (x"d0",x"49",x"e8",x"d3"),
  3175 => (x"e5",x"c0",x"81",x"66"),
  3176 => (x"f9",x"49",x"c2",x"51"),
  3177 => (x"ff",x"cb",x"87",x"ef"),
  3178 => (x"02",x"66",x"d4",x"87"),
  3179 => (x"c3",x"87",x"ca",x"c0"),
  3180 => (x"d0",x"49",x"e8",x"d3"),
  3181 => (x"e5",x"c0",x"81",x"66"),
  3182 => (x"e0",x"ff",x"c3",x"51"),
  3183 => (x"c8",x"4a",x"c0",x"4b"),
  3184 => (x"fc",x"fc",x"49",x"c0"),
  3185 => (x"ff",x"c3",x"87",x"cc"),
  3186 => (x"50",x"cb",x"48",x"e7"),
  3187 => (x"48",x"e8",x"d3",x"c3"),
  3188 => (x"70",x"80",x"66",x"d0"),
  3189 => (x"bf",x"97",x"6e",x"7e"),
  3190 => (x"c0",x"02",x"99",x"49"),
  3191 => (x"ff",x"c3",x"87",x"cc"),
  3192 => (x"50",x"c5",x"48",x"e2"),
  3193 => (x"97",x"6e",x"80",x"c9"),
  3194 => (x"1e",x"c9",x"50",x"bf"),
  3195 => (x"49",x"e0",x"ff",x"c3"),
  3196 => (x"c4",x"87",x"cc",x"f7"),
  3197 => (x"f8",x"49",x"c0",x"86"),
  3198 => (x"48",x"6e",x"87",x"db"),
  3199 => (x"e7",x"ca",x"50",x"c0"),
  3200 => (x"05",x"66",x"d4",x"87"),
  3201 => (x"d8",x"87",x"f5",x"c2"),
  3202 => (x"e8",x"c0",x"48",x"66"),
  3203 => (x"c0",x"c1",x"05",x"a8"),
  3204 => (x"49",x"66",x"dc",x"87"),
  3205 => (x"c0",x"c0",x"c0",x"c1"),
  3206 => (x"e0",x"c0",x"91",x"c0"),
  3207 => (x"c0",x"d0",x"4a",x"66"),
  3208 => (x"a1",x"72",x"92",x"c0"),
  3209 => (x"97",x"66",x"c4",x"49"),
  3210 => (x"c0",x"c4",x"4a",x"bf"),
  3211 => (x"49",x"a1",x"72",x"92"),
  3212 => (x"82",x"c5",x"4a",x"6e"),
  3213 => (x"c0",x"4a",x"6a",x"97"),
  3214 => (x"72",x"48",x"a6",x"e4"),
  3215 => (x"49",x"6e",x"78",x"a1"),
  3216 => (x"69",x"97",x"81",x"c7"),
  3217 => (x"91",x"c0",x"c4",x"49"),
  3218 => (x"82",x"c8",x"4a",x"6e"),
  3219 => (x"a1",x"4a",x"6a",x"97"),
  3220 => (x"c0",x"49",x"74",x"4c"),
  3221 => (x"c0",x"81",x"66",x"e4"),
  3222 => (x"01",x"a9",x"66",x"e8"),
  3223 => (x"c0",x"87",x"cb",x"c1"),
  3224 => (x"c9",x"49",x"66",x"e4"),
  3225 => (x"d0",x"1e",x"71",x"31"),
  3226 => (x"e4",x"fd",x"49",x"66"),
  3227 => (x"86",x"c4",x"87",x"de"),
  3228 => (x"8c",x"c1",x"49",x"74"),
  3229 => (x"c0",x"02",x"99",x"71"),
  3230 => (x"66",x"cc",x"87",x"df"),
  3231 => (x"75",x"1e",x"c0",x"4d"),
  3232 => (x"f2",x"de",x"fd",x"49"),
  3233 => (x"75",x"1e",x"c1",x"87"),
  3234 => (x"ca",x"dd",x"fd",x"49"),
  3235 => (x"74",x"86",x"c8",x"87"),
  3236 => (x"71",x"8c",x"c1",x"49"),
  3237 => (x"e4",x"ff",x"05",x"99"),
  3238 => (x"f5",x"49",x"c0",x"87"),
  3239 => (x"d3",x"c3",x"87",x"f7"),
  3240 => (x"66",x"d0",x"49",x"e8"),
  3241 => (x"c7",x"51",x"c0",x"81"),
  3242 => (x"49",x"c2",x"87",x"fe"),
  3243 => (x"c3",x"87",x"e6",x"f5"),
  3244 => (x"d0",x"49",x"e8",x"d3"),
  3245 => (x"e1",x"c0",x"81",x"66"),
  3246 => (x"87",x"ec",x"c7",x"51"),
  3247 => (x"d4",x"f5",x"49",x"c2"),
  3248 => (x"e8",x"d3",x"c3",x"87"),
  3249 => (x"81",x"66",x"d0",x"49"),
  3250 => (x"c7",x"51",x"e5",x"c0"),
  3251 => (x"66",x"d4",x"87",x"da"),
  3252 => (x"87",x"fd",x"c2",x"05"),
  3253 => (x"c0",x"48",x"66",x"d8"),
  3254 => (x"c1",x"05",x"a8",x"ea"),
  3255 => (x"66",x"dc",x"87",x"c0"),
  3256 => (x"c0",x"c0",x"c1",x"49"),
  3257 => (x"c0",x"91",x"c0",x"c0"),
  3258 => (x"d0",x"4a",x"66",x"e0"),
  3259 => (x"72",x"92",x"c0",x"c0"),
  3260 => (x"66",x"c4",x"49",x"a1"),
  3261 => (x"c4",x"4a",x"bf",x"97"),
  3262 => (x"a1",x"72",x"92",x"c0"),
  3263 => (x"c5",x"4a",x"6e",x"49"),
  3264 => (x"4a",x"6a",x"97",x"82"),
  3265 => (x"48",x"a6",x"e4",x"c0"),
  3266 => (x"6e",x"78",x"a1",x"72"),
  3267 => (x"97",x"81",x"c7",x"49"),
  3268 => (x"c0",x"c4",x"49",x"69"),
  3269 => (x"c8",x"4a",x"6e",x"91"),
  3270 => (x"4a",x"6a",x"97",x"82"),
  3271 => (x"49",x"74",x"4c",x"a1"),
  3272 => (x"81",x"66",x"e4",x"c0"),
  3273 => (x"a9",x"66",x"e8",x"c0"),
  3274 => (x"87",x"d3",x"c1",x"01"),
  3275 => (x"c0",x"02",x"9c",x"74"),
  3276 => (x"66",x"cc",x"87",x"fc"),
  3277 => (x"66",x"e4",x"c0",x"4d"),
  3278 => (x"71",x"31",x"c9",x"49"),
  3279 => (x"fd",x"49",x"75",x"1e"),
  3280 => (x"c3",x"87",x"c9",x"e1"),
  3281 => (x"f2",x"49",x"e0",x"ff"),
  3282 => (x"ff",x"c3",x"87",x"eb"),
  3283 => (x"49",x"75",x"1e",x"e0"),
  3284 => (x"87",x"f2",x"dc",x"fd"),
  3285 => (x"49",x"75",x"1e",x"c1"),
  3286 => (x"87",x"fb",x"d9",x"fd"),
  3287 => (x"e4",x"c0",x"86",x"cc"),
  3288 => (x"80",x"c1",x"48",x"66"),
  3289 => (x"58",x"a6",x"e8",x"c0"),
  3290 => (x"ff",x"05",x"8c",x"c1"),
  3291 => (x"49",x"c0",x"87",x"c7"),
  3292 => (x"c3",x"87",x"e2",x"f2"),
  3293 => (x"d0",x"49",x"e8",x"d3"),
  3294 => (x"51",x"c0",x"81",x"66"),
  3295 => (x"c2",x"87",x"e9",x"c4"),
  3296 => (x"87",x"d1",x"f2",x"49"),
  3297 => (x"49",x"e8",x"d3",x"c3"),
  3298 => (x"c0",x"81",x"66",x"d0"),
  3299 => (x"d7",x"c4",x"51",x"e1"),
  3300 => (x"f1",x"49",x"c2",x"87"),
  3301 => (x"d3",x"c3",x"87",x"ff"),
  3302 => (x"66",x"d0",x"49",x"e8"),
  3303 => (x"51",x"e5",x"c0",x"81"),
  3304 => (x"c3",x"87",x"c5",x"c4"),
  3305 => (x"c0",x"4b",x"e0",x"ff"),
  3306 => (x"49",x"c0",x"c8",x"4a"),
  3307 => (x"87",x"e2",x"f4",x"fc"),
  3308 => (x"48",x"e2",x"ff",x"c3"),
  3309 => (x"49",x"74",x"50",x"c2"),
  3310 => (x"ff",x"c3",x"89",x"c5"),
  3311 => (x"c3",x"59",x"97",x"e8"),
  3312 => (x"c3",x"48",x"f4",x"d2"),
  3313 => (x"20",x"49",x"e8",x"ff"),
  3314 => (x"c3",x"41",x"20",x"41"),
  3315 => (x"c3",x"48",x"c0",x"d3"),
  3316 => (x"20",x"49",x"f0",x"ff"),
  3317 => (x"20",x"41",x"20",x"41"),
  3318 => (x"d0",x"41",x"20",x"41"),
  3319 => (x"f0",x"c0",x"49",x"66"),
  3320 => (x"c2",x"c0",x"c4",x"81"),
  3321 => (x"d3",x"c3",x"59",x"97"),
  3322 => (x"c0",x"c4",x"48",x"d4"),
  3323 => (x"41",x"20",x"49",x"c0"),
  3324 => (x"48",x"dc",x"d3",x"c3"),
  3325 => (x"49",x"c4",x"c0",x"c4"),
  3326 => (x"41",x"20",x"41",x"20"),
  3327 => (x"c0",x"02",x"66",x"d4"),
  3328 => (x"ff",x"c3",x"87",x"c7"),
  3329 => (x"ff",x"c1",x"48",x"e0"),
  3330 => (x"c1",x"49",x"74",x"50"),
  3331 => (x"c3",x"1e",x"71",x"29"),
  3332 => (x"ee",x"49",x"e0",x"ff"),
  3333 => (x"86",x"c4",x"87",x"e9"),
  3334 => (x"f8",x"ef",x"49",x"c0"),
  3335 => (x"e8",x"d3",x"c3",x"87"),
  3336 => (x"81",x"66",x"d0",x"49"),
  3337 => (x"ff",x"c1",x"51",x"c0"),
  3338 => (x"05",x"66",x"d4",x"87"),
  3339 => (x"c3",x"87",x"d2",x"c1"),
  3340 => (x"c0",x"4b",x"e0",x"ff"),
  3341 => (x"49",x"c0",x"c8",x"4a"),
  3342 => (x"87",x"d6",x"f2",x"fc"),
  3343 => (x"48",x"e3",x"ff",x"c3"),
  3344 => (x"e8",x"c0",x"50",x"c8"),
  3345 => (x"29",x"d0",x"49",x"66"),
  3346 => (x"97",x"e9",x"ff",x"c3"),
  3347 => (x"66",x"e8",x"c0",x"59"),
  3348 => (x"c3",x"29",x"c8",x"49"),
  3349 => (x"59",x"97",x"ea",x"ff"),
  3350 => (x"c0",x"80",x"c1",x"48"),
  3351 => (x"c2",x"50",x"66",x"e8"),
  3352 => (x"49",x"74",x"50",x"80"),
  3353 => (x"1e",x"71",x"29",x"c1"),
  3354 => (x"ed",x"49",x"a0",x"f5"),
  3355 => (x"86",x"c4",x"87",x"d1"),
  3356 => (x"e0",x"ee",x"49",x"c0"),
  3357 => (x"e8",x"d3",x"c3",x"87"),
  3358 => (x"81",x"66",x"d0",x"49"),
  3359 => (x"e7",x"c0",x"51",x"c0"),
  3360 => (x"e8",x"d3",x"c3",x"87"),
  3361 => (x"81",x"66",x"d0",x"49"),
  3362 => (x"c2",x"51",x"e5",x"c0"),
  3363 => (x"87",x"c5",x"ee",x"49"),
  3364 => (x"c3",x"87",x"d5",x"c0"),
  3365 => (x"d0",x"49",x"e8",x"d3"),
  3366 => (x"e0",x"c0",x"81",x"66"),
  3367 => (x"ed",x"49",x"c2",x"51"),
  3368 => (x"c3",x"c0",x"87",x"f3"),
  3369 => (x"87",x"c6",x"ee",x"87"),
  3370 => (x"26",x"8e",x"d4",x"ff"),
  3371 => (x"26",x"4c",x"26",x"4d"),
  3372 => (x"00",x"4f",x"26",x"4b"),
  3373 => (x"34",x"36",x"43",x"54"),
  3374 => (x"20",x"20",x"20",x"20"),
  3375 => (x"00",x"00",x"00",x"00"),
  3376 => (x"69",x"4d",x"65",x"44"),
  3377 => (x"66",x"69",x"54",x"53"),
  3378 => (x"44",x"48",x"20",x"79"),
  3379 => (x"20",x"30",x"20",x"44"),
  3380 => (x"00",x"00",x"00",x"00"),
  3381 => (x"20",x"32",x"33",x"38"),
  3382 => (x"00",x"00",x"00",x"00"),
  3383 => (x"32",x"31",x"30",x"32"),
  3384 => (x"39",x"32",x"39",x"30"),
  3385 => (x"00",x"00",x"00",x"09"),
  3386 => (x"73",x"1e",x"00",x"00"),
  3387 => (x"ff",x"86",x"e0",x"1e"),
  3388 => (x"c5",x"c8",x"48",x"d0"),
  3389 => (x"48",x"d4",x"ff",x"78"),
  3390 => (x"1e",x"d0",x"78",x"c5"),
  3391 => (x"49",x"4b",x"a6",x"c4"),
  3392 => (x"87",x"e3",x"f1",x"fc"),
  3393 => (x"d0",x"ff",x"86",x"c4"),
  3394 => (x"ca",x"78",x"c4",x"48"),
  3395 => (x"c1",x"49",x"66",x"97"),
  3396 => (x"87",x"c5",x"02",x"99"),
  3397 => (x"e8",x"ec",x"49",x"73"),
  3398 => (x"26",x"8e",x"e0",x"87"),
  3399 => (x"1e",x"4f",x"26",x"4b"),
  3400 => (x"c4",x"4a",x"d4",x"ff"),
  3401 => (x"c4",x"48",x"c8",x"d8"),
  3402 => (x"78",x"bf",x"f4",x"d1"),
  3403 => (x"ff",x"7a",x"ff",x"c3"),
  3404 => (x"78",x"c5",x"48",x"d0"),
  3405 => (x"d1",x"c4",x"7a",x"c4"),
  3406 => (x"48",x"49",x"bf",x"f4"),
  3407 => (x"7a",x"70",x"28",x"d8"),
  3408 => (x"28",x"d0",x"48",x"71"),
  3409 => (x"48",x"71",x"7a",x"70"),
  3410 => (x"7a",x"70",x"28",x"c8"),
  3411 => (x"bf",x"f4",x"d1",x"c4"),
  3412 => (x"48",x"d0",x"ff",x"7a"),
  3413 => (x"4f",x"26",x"78",x"c4"),
  3414 => (x"c4",x"4a",x"c0",x"1e"),
  3415 => (x"02",x"bf",x"fc",x"d8"),
  3416 => (x"c4",x"49",x"87",x"ca"),
  3417 => (x"c1",x"48",x"fc",x"d8"),
  3418 => (x"4a",x"11",x"78",x"a1"),
  3419 => (x"c6",x"05",x"9a",x"72"),
  3420 => (x"fc",x"d8",x"c4",x"87"),
  3421 => (x"72",x"78",x"c0",x"48"),
  3422 => (x"1e",x"4f",x"26",x"48"),
  3423 => (x"48",x"fc",x"d8",x"c4"),
  3424 => (x"bf",x"d8",x"f4",x"c3"),
  3425 => (x"0e",x"4f",x"26",x"78"),
  3426 => (x"0e",x"5c",x"5b",x"5e"),
  3427 => (x"d0",x"ff",x"4a",x"71"),
  3428 => (x"4b",x"d4",x"ff",x"4c"),
  3429 => (x"d5",x"c1",x"7c",x"c5"),
  3430 => (x"7b",x"66",x"cc",x"7b"),
  3431 => (x"7c",x"c5",x"7c",x"c4"),
  3432 => (x"c1",x"7b",x"d3",x"c1"),
  3433 => (x"c8",x"7c",x"c4",x"7b"),
  3434 => (x"d4",x"c1",x"7c",x"c5"),
  3435 => (x"b7",x"49",x"c0",x"7b"),
  3436 => (x"87",x"ca",x"06",x"aa"),
  3437 => (x"81",x"c1",x"7b",x"c0"),
  3438 => (x"04",x"a9",x"b7",x"72"),
  3439 => (x"7c",x"c4",x"87",x"f6"),
  3440 => (x"d3",x"c1",x"7c",x"c5"),
  3441 => (x"c4",x"7b",x"c0",x"7b"),
  3442 => (x"26",x"4c",x"26",x"7c"),
  3443 => (x"1e",x"4f",x"26",x"4b"),
  3444 => (x"4b",x"71",x"1e",x"73"),
  3445 => (x"97",x"e0",x"f3",x"c1"),
  3446 => (x"b7",x"c2",x"49",x"bf"),
  3447 => (x"f3",x"c0",x"03",x"a9"),
  3448 => (x"c4",x"1e",x"73",x"87"),
  3449 => (x"fd",x"49",x"dc",x"cc"),
  3450 => (x"c4",x"87",x"c8",x"cb"),
  3451 => (x"02",x"98",x"70",x"86"),
  3452 => (x"c4",x"87",x"e1",x"c0"),
  3453 => (x"4a",x"bf",x"e4",x"cc"),
  3454 => (x"c0",x"c3",x"2a",x"ca"),
  3455 => (x"87",x"ce",x"02",x"8a"),
  3456 => (x"05",x"8a",x"c0",x"c1"),
  3457 => (x"f3",x"c1",x"87",x"ce"),
  3458 => (x"50",x"c0",x"48",x"e0"),
  3459 => (x"f3",x"c1",x"87",x"c6"),
  3460 => (x"50",x"c1",x"48",x"e0"),
  3461 => (x"4f",x"26",x"4b",x"26"),
  3462 => (x"71",x"1e",x"73",x"1e"),
  3463 => (x"c6",x"02",x"9a",x"4a"),
  3464 => (x"cc",x"dd",x"c3",x"87"),
  3465 => (x"c3",x"78",x"c0",x"48"),
  3466 => (x"49",x"bf",x"c8",x"dd"),
  3467 => (x"87",x"c0",x"ce",x"ff"),
  3468 => (x"c4",x"02",x"98",x"70"),
  3469 => (x"49",x"d4",x"87",x"cd"),
  3470 => (x"87",x"e8",x"cd",x"ff"),
  3471 => (x"58",x"cc",x"dd",x"c3"),
  3472 => (x"bf",x"cc",x"dd",x"c3"),
  3473 => (x"87",x"fb",x"c0",x"05"),
  3474 => (x"49",x"e0",x"d1",x"c4"),
  3475 => (x"87",x"cb",x"df",x"fe"),
  3476 => (x"04",x"a8",x"b7",x"c0"),
  3477 => (x"d1",x"c4",x"87",x"ce"),
  3478 => (x"de",x"fe",x"49",x"e0"),
  3479 => (x"b7",x"c0",x"87",x"fd"),
  3480 => (x"87",x"f2",x"03",x"a8"),
  3481 => (x"bf",x"cc",x"dd",x"c3"),
  3482 => (x"cc",x"dd",x"c3",x"49"),
  3483 => (x"78",x"a1",x"c1",x"48"),
  3484 => (x"81",x"dc",x"f4",x"c3"),
  3485 => (x"dd",x"c3",x"48",x"11"),
  3486 => (x"dd",x"c3",x"58",x"d4"),
  3487 => (x"78",x"c0",x"48",x"d4"),
  3488 => (x"c3",x"87",x"c0",x"c3"),
  3489 => (x"02",x"bf",x"d4",x"dd"),
  3490 => (x"c4",x"87",x"f5",x"c1"),
  3491 => (x"fe",x"49",x"e0",x"d1"),
  3492 => (x"c0",x"87",x"c8",x"de"),
  3493 => (x"cd",x"04",x"a8",x"b7"),
  3494 => (x"d4",x"dd",x"c3",x"87"),
  3495 => (x"88",x"c1",x"48",x"bf"),
  3496 => (x"58",x"d8",x"dd",x"c3"),
  3497 => (x"d7",x"c4",x"87",x"dd"),
  3498 => (x"ff",x"49",x"bf",x"c0"),
  3499 => (x"70",x"87",x"c1",x"cc"),
  3500 => (x"ce",x"c0",x"02",x"98"),
  3501 => (x"e0",x"d1",x"c4",x"87"),
  3502 => (x"d3",x"db",x"fe",x"49"),
  3503 => (x"cc",x"dd",x"c3",x"87"),
  3504 => (x"c3",x"78",x"c0",x"48"),
  3505 => (x"05",x"bf",x"d0",x"dd"),
  3506 => (x"c3",x"87",x"f8",x"c1"),
  3507 => (x"05",x"bf",x"d4",x"dd"),
  3508 => (x"c3",x"87",x"f0",x"c1"),
  3509 => (x"49",x"bf",x"cc",x"dd"),
  3510 => (x"48",x"cc",x"dd",x"c3"),
  3511 => (x"c3",x"78",x"a1",x"c1"),
  3512 => (x"11",x"81",x"dc",x"f4"),
  3513 => (x"c0",x"c2",x"49",x"4b"),
  3514 => (x"cc",x"c0",x"02",x"99"),
  3515 => (x"c1",x"48",x"73",x"87"),
  3516 => (x"dd",x"c3",x"98",x"ff"),
  3517 => (x"ca",x"c1",x"58",x"d8"),
  3518 => (x"d4",x"dd",x"c3",x"87"),
  3519 => (x"87",x"c3",x"c1",x"5b"),
  3520 => (x"bf",x"d0",x"dd",x"c3"),
  3521 => (x"87",x"fb",x"c0",x"02"),
  3522 => (x"bf",x"cc",x"dd",x"c3"),
  3523 => (x"cc",x"dd",x"c3",x"49"),
  3524 => (x"78",x"a1",x"c1",x"48"),
  3525 => (x"81",x"dc",x"f4",x"c3"),
  3526 => (x"1e",x"49",x"69",x"97"),
  3527 => (x"49",x"e0",x"d1",x"c4"),
  3528 => (x"87",x"c3",x"da",x"fe"),
  3529 => (x"dd",x"c3",x"86",x"c4"),
  3530 => (x"c1",x"48",x"bf",x"d0"),
  3531 => (x"d4",x"dd",x"c3",x"88"),
  3532 => (x"d4",x"dd",x"c3",x"58"),
  3533 => (x"c0",x"78",x"c1",x"48"),
  3534 => (x"ff",x"49",x"ec",x"f6"),
  3535 => (x"c4",x"87",x"e5",x"c9"),
  3536 => (x"26",x"58",x"c4",x"d7"),
  3537 => (x"00",x"4f",x"26",x"4b"),
  3538 => (x"00",x"00",x"00",x"00"),
  3539 => (x"00",x"00",x"00",x"00"),
  3540 => (x"00",x"00",x"00",x"00"),
  3541 => (x"00",x"00",x"00",x"00"),
  3542 => (x"71",x"1e",x"73",x"1e"),
  3543 => (x"fb",x"fd",x"49",x"4b"),
  3544 => (x"d2",x"c4",x"87",x"e8"),
  3545 => (x"02",x"bf",x"97",x"c8"),
  3546 => (x"1e",x"c3",x"87",x"cb"),
  3547 => (x"49",x"c0",x"c0",x"c4"),
  3548 => (x"c4",x"87",x"d4",x"f8"),
  3549 => (x"fd",x"49",x"73",x"86"),
  3550 => (x"26",x"87",x"cf",x"fb"),
  3551 => (x"1e",x"4f",x"26",x"4b"),
  3552 => (x"da",x"f6",x"1e",x"73"),
  3553 => (x"49",x"f4",x"c7",x"87"),
  3554 => (x"87",x"d8",x"c8",x"ff"),
  3555 => (x"ff",x"49",x"4b",x"70"),
  3556 => (x"70",x"87",x"dd",x"c8"),
  3557 => (x"87",x"cb",x"05",x"98"),
  3558 => (x"c8",x"ff",x"49",x"73"),
  3559 => (x"98",x"70",x"87",x"d2"),
  3560 => (x"26",x"87",x"f5",x"02"),
  3561 => (x"0e",x"4f",x"26",x"4b"),
  3562 => (x"5d",x"5c",x"5b",x"5e"),
  3563 => (x"71",x"86",x"f8",x"0e"),
  3564 => (x"fd",x"4d",x"c0",x"4b"),
  3565 => (x"70",x"87",x"e7",x"d4"),
  3566 => (x"02",x"9b",x"73",x"4c"),
  3567 => (x"c1",x"87",x"c2",x"c5"),
  3568 => (x"c1",x"48",x"e0",x"f3"),
  3569 => (x"c4",x"1e",x"73",x"50"),
  3570 => (x"fd",x"49",x"dc",x"cc"),
  3571 => (x"c4",x"87",x"e4",x"c3"),
  3572 => (x"02",x"98",x"70",x"86"),
  3573 => (x"c4",x"87",x"ff",x"c3"),
  3574 => (x"48",x"bf",x"f4",x"d1"),
  3575 => (x"d1",x"c4",x"b0",x"c1"),
  3576 => (x"fa",x"f4",x"58",x"f8"),
  3577 => (x"e0",x"ff",x"c3",x"87"),
  3578 => (x"dc",x"cc",x"c4",x"1e"),
  3579 => (x"c6",x"c9",x"fd",x"49"),
  3580 => (x"c3",x"86",x"c4",x"87"),
  3581 => (x"7e",x"bf",x"ec",x"ff"),
  3582 => (x"c3",x"48",x"a6",x"c4"),
  3583 => (x"78",x"bf",x"f0",x"ff"),
  3584 => (x"97",x"e0",x"ff",x"c3"),
  3585 => (x"a9",x"c1",x"49",x"bf"),
  3586 => (x"87",x"ca",x"c3",x"05"),
  3587 => (x"bf",x"e4",x"ff",x"c3"),
  3588 => (x"71",x"b1",x"c1",x"49"),
  3589 => (x"ff",x"cf",x"ff",x"48"),
  3590 => (x"f8",x"d1",x"c4",x"98"),
  3591 => (x"e1",x"ff",x"c3",x"58"),
  3592 => (x"c2",x"48",x"bf",x"97"),
  3593 => (x"c3",x"58",x"d8",x"e6"),
  3594 => (x"49",x"bf",x"e8",x"ff"),
  3595 => (x"87",x"ef",x"dd",x"fd"),
  3596 => (x"c0",x"02",x"98",x"70"),
  3597 => (x"ff",x"c3",x"87",x"e2"),
  3598 => (x"cc",x"c4",x"1e",x"e0"),
  3599 => (x"c7",x"fd",x"49",x"dc"),
  3600 => (x"ff",x"c3",x"87",x"f5"),
  3601 => (x"fd",x"49",x"bf",x"e8"),
  3602 => (x"c0",x"87",x"f4",x"d0"),
  3603 => (x"f4",x"ff",x"c3",x"1e"),
  3604 => (x"87",x"cc",x"c4",x"49"),
  3605 => (x"4d",x"70",x"86",x"c8"),
  3606 => (x"d0",x"fd",x"49",x"74"),
  3607 => (x"1e",x"73",x"87",x"e1"),
  3608 => (x"49",x"dc",x"cc",x"c4"),
  3609 => (x"87",x"cb",x"c1",x"fd"),
  3610 => (x"49",x"6e",x"86",x"c4"),
  3611 => (x"87",x"ef",x"dc",x"fd"),
  3612 => (x"c0",x"02",x"98",x"70"),
  3613 => (x"ff",x"c3",x"87",x"e1"),
  3614 => (x"cc",x"c4",x"1e",x"e0"),
  3615 => (x"c6",x"fd",x"49",x"dc"),
  3616 => (x"ff",x"c3",x"87",x"f5"),
  3617 => (x"fd",x"49",x"bf",x"ec"),
  3618 => (x"c0",x"87",x"f4",x"cf"),
  3619 => (x"c0",x"c4",x"1e",x"f2"),
  3620 => (x"cb",x"c3",x"49",x"c0"),
  3621 => (x"74",x"86",x"c8",x"87"),
  3622 => (x"e2",x"cf",x"fd",x"49"),
  3623 => (x"c4",x"1e",x"73",x"87"),
  3624 => (x"fd",x"49",x"dc",x"cc"),
  3625 => (x"c4",x"87",x"cc",x"c0"),
  3626 => (x"fd",x"49",x"66",x"86"),
  3627 => (x"70",x"87",x"f0",x"db"),
  3628 => (x"e1",x"c0",x"02",x"98"),
  3629 => (x"e0",x"ff",x"c3",x"87"),
  3630 => (x"dc",x"cc",x"c4",x"1e"),
  3631 => (x"f6",x"c5",x"fd",x"49"),
  3632 => (x"f0",x"ff",x"c3",x"87"),
  3633 => (x"ce",x"fd",x"49",x"bf"),
  3634 => (x"f3",x"c0",x"87",x"f5"),
  3635 => (x"cc",x"c0",x"c4",x"1e"),
  3636 => (x"87",x"cc",x"c2",x"49"),
  3637 => (x"1e",x"c2",x"86",x"c8"),
  3638 => (x"49",x"c0",x"c0",x"c4"),
  3639 => (x"c3",x"87",x"e8",x"f2"),
  3640 => (x"c0",x"c0",x"c4",x"1e"),
  3641 => (x"87",x"df",x"f2",x"49"),
  3642 => (x"d1",x"c4",x"86",x"c8"),
  3643 => (x"fe",x"48",x"bf",x"f4"),
  3644 => (x"f8",x"d1",x"c4",x"98"),
  3645 => (x"87",x"e7",x"f0",x"58"),
  3646 => (x"bf",x"d4",x"e6",x"c2"),
  3647 => (x"d2",x"f5",x"fe",x"49"),
  3648 => (x"f8",x"48",x"75",x"87"),
  3649 => (x"26",x"4d",x"26",x"8e"),
  3650 => (x"26",x"4b",x"26",x"4c"),
  3651 => (x"1e",x"73",x"1e",x"4f"),
  3652 => (x"49",x"ca",x"4b",x"71"),
  3653 => (x"87",x"f6",x"dc",x"fc"),
  3654 => (x"cc",x"c4",x"1e",x"73"),
  3655 => (x"fe",x"fc",x"49",x"dc"),
  3656 => (x"86",x"c4",x"87",x"d1"),
  3657 => (x"c0",x"02",x"98",x"70"),
  3658 => (x"d8",x"c4",x"87",x"f0"),
  3659 => (x"50",x"c1",x"48",x"c4"),
  3660 => (x"bf",x"d4",x"e6",x"c2"),
  3661 => (x"c4",x"80",x"c2",x"50"),
  3662 => (x"78",x"bf",x"f4",x"d1"),
  3663 => (x"50",x"c0",x"80",x"db"),
  3664 => (x"50",x"c0",x"80",x"cb"),
  3665 => (x"50",x"c0",x"80",x"cb"),
  3666 => (x"1e",x"a0",x"c8",x"ff"),
  3667 => (x"49",x"dc",x"cc",x"c4"),
  3668 => (x"87",x"f2",x"c4",x"fd"),
  3669 => (x"48",x"c1",x"86",x"c4"),
  3670 => (x"48",x"c0",x"87",x"c2"),
  3671 => (x"4f",x"26",x"4b",x"26"),
  3672 => (x"5c",x"5b",x"5e",x"0e"),
  3673 => (x"86",x"f4",x"0e",x"5d"),
  3674 => (x"a6",x"c4",x"7e",x"71"),
  3675 => (x"dc",x"78",x"c0",x"48"),
  3676 => (x"f0",x"c0",x"4d",x"66"),
  3677 => (x"02",x"66",x"dc",x"8d"),
  3678 => (x"75",x"87",x"e6",x"c0"),
  3679 => (x"f6",x"c1",x"02",x"9d"),
  3680 => (x"8c",x"c1",x"4c",x"87"),
  3681 => (x"87",x"ef",x"c1",x"02"),
  3682 => (x"d5",x"c2",x"02",x"8c"),
  3683 => (x"c2",x"02",x"8c",x"87"),
  3684 => (x"8c",x"d0",x"87",x"d0"),
  3685 => (x"87",x"eb",x"c4",x"02"),
  3686 => (x"c4",x"02",x"8c",x"c1"),
  3687 => (x"f5",x"c4",x"87",x"f0"),
  3688 => (x"c4",x"02",x"6e",x"87"),
  3689 => (x"97",x"6e",x"87",x"f0"),
  3690 => (x"e9",x"c4",x"02",x"bf"),
  3691 => (x"c4",x"1e",x"c2",x"87"),
  3692 => (x"ef",x"49",x"c0",x"c0"),
  3693 => (x"86",x"c4",x"87",x"d1"),
  3694 => (x"4b",x"d8",x"d8",x"c4"),
  3695 => (x"49",x"cb",x"4a",x"6e"),
  3696 => (x"87",x"fe",x"db",x"fc"),
  3697 => (x"48",x"e3",x"d8",x"c4"),
  3698 => (x"cc",x"fd",x"50",x"c0"),
  3699 => (x"d8",x"c4",x"87",x"d0"),
  3700 => (x"d1",x"c4",x"58",x"d0"),
  3701 => (x"c1",x"48",x"bf",x"f4"),
  3702 => (x"f8",x"d1",x"c4",x"b0"),
  3703 => (x"87",x"ff",x"ec",x"58"),
  3704 => (x"49",x"d8",x"d8",x"c4"),
  3705 => (x"c4",x"87",x"e8",x"ef"),
  3706 => (x"fd",x"49",x"d8",x"d8"),
  3707 => (x"c4",x"87",x"d6",x"e0"),
  3708 => (x"78",x"c1",x"48",x"a6"),
  3709 => (x"75",x"87",x"df",x"c3"),
  3710 => (x"ff",x"49",x"c0",x"1e"),
  3711 => (x"75",x"87",x"d5",x"c4"),
  3712 => (x"87",x"fb",x"f5",x"49"),
  3713 => (x"66",x"c8",x"1e",x"75"),
  3714 => (x"c7",x"c4",x"ff",x"49"),
  3715 => (x"75",x"86",x"c8",x"87"),
  3716 => (x"91",x"c8",x"c1",x"49"),
  3717 => (x"81",x"e0",x"d2",x"c4"),
  3718 => (x"a6",x"c4",x"81",x"c8"),
  3719 => (x"c2",x"78",x"69",x"48"),
  3720 => (x"49",x"75",x"87",x"f4"),
  3721 => (x"c4",x"91",x"c8",x"c1"),
  3722 => (x"71",x"48",x"e0",x"d2"),
  3723 => (x"58",x"a6",x"c8",x"80"),
  3724 => (x"c8",x"48",x"66",x"c4"),
  3725 => (x"58",x"a6",x"cc",x"80"),
  3726 => (x"c0",x"48",x"66",x"c8"),
  3727 => (x"c0",x"02",x"6e",x"78"),
  3728 => (x"4c",x"75",x"87",x"e5"),
  3729 => (x"d8",x"c4",x"94",x"cc"),
  3730 => (x"4b",x"74",x"84",x"cc"),
  3731 => (x"49",x"cb",x"4a",x"6e"),
  3732 => (x"87",x"ee",x"d9",x"fc"),
  3733 => (x"c0",x"49",x"a4",x"cb"),
  3734 => (x"c8",x"1e",x"74",x"51"),
  3735 => (x"f9",x"fc",x"49",x"66"),
  3736 => (x"86",x"c4",x"87",x"d1"),
  3737 => (x"75",x"87",x"ca",x"c0"),
  3738 => (x"c4",x"91",x"cc",x"49"),
  3739 => (x"c0",x"81",x"cc",x"d8"),
  3740 => (x"e9",x"c9",x"fd",x"51"),
  3741 => (x"75",x"4a",x"70",x"87"),
  3742 => (x"c4",x"91",x"c4",x"49"),
  3743 => (x"72",x"81",x"c8",x"d8"),
  3744 => (x"bf",x"66",x"c8",x"79"),
  3745 => (x"87",x"d9",x"c0",x"02"),
  3746 => (x"89",x"c2",x"49",x"75"),
  3747 => (x"71",x"48",x"c0",x"d0"),
  3748 => (x"c4",x"49",x"70",x"30"),
  3749 => (x"48",x"bf",x"f4",x"d1"),
  3750 => (x"d1",x"c4",x"b0",x"71"),
  3751 => (x"d8",x"c0",x"58",x"f8"),
  3752 => (x"c2",x"49",x"75",x"87"),
  3753 => (x"48",x"c0",x"d0",x"89"),
  3754 => (x"49",x"70",x"30",x"71"),
  3755 => (x"d1",x"c4",x"b9",x"ff"),
  3756 => (x"71",x"48",x"bf",x"f4"),
  3757 => (x"f8",x"d1",x"c4",x"98"),
  3758 => (x"48",x"a6",x"c4",x"58"),
  3759 => (x"78",x"bf",x"66",x"c8"),
  3760 => (x"6e",x"87",x"d3",x"c0"),
  3761 => (x"87",x"df",x"f3",x"49"),
  3762 => (x"c0",x"58",x"a6",x"c8"),
  3763 => (x"49",x"6e",x"87",x"c8"),
  3764 => (x"c8",x"87",x"fa",x"f8"),
  3765 => (x"d1",x"c4",x"58",x"a6"),
  3766 => (x"fe",x"48",x"bf",x"f4"),
  3767 => (x"f8",x"d1",x"c4",x"98"),
  3768 => (x"87",x"fb",x"e8",x"58"),
  3769 => (x"f4",x"48",x"66",x"c4"),
  3770 => (x"26",x"4d",x"26",x"8e"),
  3771 => (x"26",x"4b",x"26",x"4c"),
  3772 => (x"1e",x"73",x"1e",x"4f"),
  3773 => (x"48",x"f4",x"d1",x"c4"),
  3774 => (x"f3",x"c1",x"78",x"c1"),
  3775 => (x"50",x"c1",x"48",x"e0"),
  3776 => (x"48",x"c4",x"c8",x"c1"),
  3777 => (x"d6",x"e8",x"50",x"c0"),
  3778 => (x"c4",x"1e",x"c3",x"87"),
  3779 => (x"e9",x"49",x"c0",x"c0"),
  3780 => (x"1e",x"c2",x"87",x"f5"),
  3781 => (x"49",x"c0",x"c0",x"c4"),
  3782 => (x"c8",x"87",x"ec",x"e9"),
  3783 => (x"f0",x"f4",x"c3",x"86"),
  3784 => (x"c2",x"f2",x"49",x"bf"),
  3785 => (x"05",x"98",x"70",x"87"),
  3786 => (x"e7",x"87",x"ef",x"c1"),
  3787 => (x"f4",x"c3",x"87",x"f1"),
  3788 => (x"ea",x"49",x"bf",x"ec"),
  3789 => (x"f4",x"c3",x"87",x"d9"),
  3790 => (x"fd",x"49",x"bf",x"ec"),
  3791 => (x"c4",x"87",x"c6",x"db"),
  3792 => (x"48",x"bf",x"f4",x"d1"),
  3793 => (x"d1",x"c4",x"98",x"fe"),
  3794 => (x"d2",x"e7",x"58",x"f8"),
  3795 => (x"49",x"d0",x"c6",x"87"),
  3796 => (x"87",x"d0",x"f9",x"fe"),
  3797 => (x"fe",x"49",x"4b",x"70"),
  3798 => (x"70",x"87",x"d5",x"f9"),
  3799 => (x"87",x"cc",x"05",x"98"),
  3800 => (x"f9",x"fe",x"49",x"73"),
  3801 => (x"98",x"70",x"87",x"ca"),
  3802 => (x"87",x"f4",x"ff",x"02"),
  3803 => (x"bf",x"f4",x"d1",x"c4"),
  3804 => (x"c4",x"b0",x"c1",x"48"),
  3805 => (x"e6",x"58",x"f8",x"d1"),
  3806 => (x"e4",x"c1",x"87",x"e5"),
  3807 => (x"e3",x"f8",x"fe",x"49"),
  3808 => (x"49",x"4b",x"70",x"87"),
  3809 => (x"87",x"e8",x"f8",x"fe"),
  3810 => (x"c0",x"05",x"98",x"70"),
  3811 => (x"49",x"73",x"87",x"cc"),
  3812 => (x"87",x"dc",x"f8",x"fe"),
  3813 => (x"ff",x"02",x"98",x"70"),
  3814 => (x"d1",x"c4",x"87",x"f4"),
  3815 => (x"fe",x"48",x"bf",x"f4"),
  3816 => (x"f8",x"d1",x"c4",x"98"),
  3817 => (x"87",x"f7",x"e5",x"58"),
  3818 => (x"87",x"f4",x"cf",x"ff"),
  3819 => (x"87",x"d0",x"c7",x"fe"),
  3820 => (x"e3",x"e9",x"49",x"c1"),
  3821 => (x"26",x"48",x"c0",x"87"),
  3822 => (x"1e",x"4f",x"26",x"4b"),
  3823 => (x"4b",x"71",x"1e",x"73"),
  3824 => (x"87",x"c8",x"c4",x"ff"),
  3825 => (x"cf",x"fe",x"49",x"73"),
  3826 => (x"4b",x"26",x"87",x"c6"),
  3827 => (x"5e",x"0e",x"4f",x"26"),
  3828 => (x"fc",x"0e",x"5c",x"5b"),
  3829 => (x"ff",x"ff",x"c1",x"86"),
  3830 => (x"c0",x"4b",x"6e",x"4c"),
  3831 => (x"87",x"f8",x"e8",x"49"),
  3832 => (x"87",x"d7",x"ed",x"fe"),
  3833 => (x"87",x"d5",x"f9",x"fe"),
  3834 => (x"73",x"87",x"ff",x"e3"),
  3835 => (x"c1",x"99",x"74",x"49"),
  3836 => (x"05",x"99",x"71",x"83"),
  3837 => (x"ff",x"fd",x"87",x"e5"),
  3838 => (x"49",x"70",x"87",x"ea"),
  3839 => (x"87",x"e7",x"d4",x"fe"),
  3840 => (x"fc",x"87",x"d8",x"ff"),
  3841 => (x"26",x"4c",x"26",x"8e"),
  3842 => (x"00",x"4f",x"26",x"4b"),
  3843 => (x"f5",x"f2",x"eb",x"f4"),
  3844 => (x"0c",x"04",x"06",x"05"),
  3845 => (x"0a",x"83",x"0b",x"03"),
  3846 => (x"00",x"00",x"00",x"66"),
  3847 => (x"00",x"da",x"00",x"5a"),
  3848 => (x"08",x"94",x"80",x"00"),
  3849 => (x"00",x"78",x"80",x"05"),
  3850 => (x"00",x"01",x"80",x"02"),
  3851 => (x"00",x"09",x"80",x"03"),
  3852 => (x"00",x"00",x"80",x"04"),
  3853 => (x"08",x"91",x"80",x"01"),
  3854 => (x"00",x"00",x"00",x"26"),
  3855 => (x"00",x"00",x"00",x"1d"),
  3856 => (x"00",x"00",x"00",x"1c"),
  3857 => (x"00",x"00",x"00",x"25"),
  3858 => (x"00",x"00",x"00",x"1a"),
  3859 => (x"00",x"00",x"00",x"1b"),
  3860 => (x"00",x"00",x"00",x"24"),
  3861 => (x"00",x"00",x"01",x"12"),
  3862 => (x"00",x"00",x"00",x"2e"),
  3863 => (x"00",x"00",x"00",x"2d"),
  3864 => (x"00",x"00",x"00",x"23"),
  3865 => (x"00",x"00",x"00",x"36"),
  3866 => (x"00",x"00",x"00",x"21"),
  3867 => (x"00",x"00",x"00",x"2b"),
  3868 => (x"00",x"00",x"00",x"2c"),
  3869 => (x"00",x"00",x"00",x"22"),
  3870 => (x"00",x"6c",x"00",x"3d"),
  3871 => (x"00",x"00",x"00",x"35"),
  3872 => (x"00",x"00",x"00",x"34"),
  3873 => (x"00",x"75",x"00",x"3e"),
  3874 => (x"00",x"00",x"00",x"32"),
  3875 => (x"00",x"00",x"00",x"33"),
  3876 => (x"00",x"6b",x"00",x"3c"),
  3877 => (x"00",x"00",x"00",x"2a"),
  3878 => (x"00",x"7d",x"00",x"46"),
  3879 => (x"00",x"73",x"00",x"43"),
  3880 => (x"00",x"69",x"00",x"3b"),
  3881 => (x"00",x"ca",x"00",x"45"),
  3882 => (x"00",x"70",x"00",x"3a"),
  3883 => (x"00",x"72",x"00",x"42"),
  3884 => (x"00",x"74",x"00",x"44"),
  3885 => (x"00",x"00",x"00",x"31"),
  3886 => (x"00",x"00",x"00",x"55"),
  3887 => (x"00",x"7c",x"00",x"4d"),
  3888 => (x"00",x"7a",x"00",x"4b"),
  3889 => (x"00",x"00",x"00",x"7b"),
  3890 => (x"00",x"71",x"00",x"49"),
  3891 => (x"00",x"84",x"00",x"4c"),
  3892 => (x"00",x"77",x"00",x"54"),
  3893 => (x"00",x"00",x"00",x"41"),
  3894 => (x"00",x"00",x"00",x"61"),
  3895 => (x"00",x"7c",x"00",x"5b"),
  3896 => (x"00",x"00",x"00",x"52"),
  3897 => (x"00",x"00",x"00",x"f1"),
  3898 => (x"00",x"00",x"02",x"59"),
  3899 => (x"00",x"5d",x"00",x"0e"),
  3900 => (x"00",x"00",x"00",x"5d"),
  3901 => (x"00",x"79",x"00",x"4a"),
  3902 => (x"00",x"00",x"00",x"16"),
  3903 => (x"00",x"07",x"00",x"76"),
  3904 => (x"00",x"0d",x"04",x"14"),
  3905 => (x"00",x"00",x"00",x"1e"),
  3906 => (x"00",x"00",x"00",x"29"),
  3907 => (x"00",x"00",x"00",x"11"),
  3908 => (x"00",x"00",x"00",x"15"),
  3909 => (x"00",x"00",x"40",x"00"),
  3910 => (x"00",x"00",x"3d",x"34"),
  3911 => (x"08",x"82",x"ff",x"01"),
  3912 => (x"64",x"f3",x"c8",x"f3"),
  3913 => (x"01",x"f2",x"50",x"f3"),
  3914 => (x"00",x"f4",x"01",x"81"),
  3915 => (x"00",x"00",x"3f",x"a0"),
  3916 => (x"00",x"00",x"3f",x"ac"),
  3917 => (x"72",x"61",x"74",x"41"),
  3918 => (x"54",x"53",x"20",x"69"),
  3919 => (x"31",x"50",x"3b",x"3b"),
  3920 => (x"6f",x"74",x"53",x"2c"),
  3921 => (x"65",x"67",x"61",x"72"),
  3922 => (x"53",x"31",x"50",x"3b"),
  3923 => (x"53",x"2c",x"55",x"30"),
  3924 => (x"46",x"2c",x"20",x"54"),
  3925 => (x"70",x"70",x"6f",x"6c"),
  3926 => (x"3a",x"41",x"20",x"79"),
  3927 => (x"53",x"31",x"50",x"3b"),
  3928 => (x"53",x"2c",x"55",x"31"),
  3929 => (x"46",x"2c",x"20",x"54"),
  3930 => (x"70",x"70",x"6f",x"6c"),
  3931 => (x"3a",x"42",x"20",x"79"),
  3932 => (x"4f",x"31",x"50",x"3b"),
  3933 => (x"57",x"2c",x"37",x"36"),
  3934 => (x"65",x"74",x"69",x"72"),
  3935 => (x"6f",x"72",x"70",x"20"),
  3936 => (x"74",x"63",x"65",x"74"),
  3937 => (x"66",x"66",x"4f",x"2c"),
  3938 => (x"2c",x"3a",x"41",x"2c"),
  3939 => (x"42",x"2c",x"3a",x"42"),
  3940 => (x"3b",x"68",x"74",x"6f"),
  3941 => (x"41",x"4f",x"31",x"50"),
  3942 => (x"61",x"48",x"2c",x"42"),
  3943 => (x"64",x"20",x"64",x"72"),
  3944 => (x"73",x"6b",x"73",x"69"),
  3945 => (x"6e",x"6f",x"4e",x"2c"),
  3946 => (x"6e",x"55",x"2c",x"65"),
  3947 => (x"30",x"20",x"74",x"69"),
  3948 => (x"69",x"6e",x"55",x"2c"),
  3949 => (x"2c",x"31",x"20",x"74"),
  3950 => (x"68",x"74",x"6f",x"42"),
  3951 => (x"53",x"31",x"50",x"3b"),
  3952 => (x"48",x"2c",x"55",x"32"),
  3953 => (x"48",x"56",x"46",x"44"),
  3954 => (x"61",x"48",x"2c",x"44"),
  3955 => (x"69",x"66",x"64",x"72"),
  3956 => (x"30",x"20",x"65",x"6c"),
  3957 => (x"53",x"31",x"50",x"3b"),
  3958 => (x"48",x"2c",x"55",x"33"),
  3959 => (x"48",x"56",x"46",x"44"),
  3960 => (x"61",x"48",x"2c",x"44"),
  3961 => (x"69",x"66",x"64",x"72"),
  3962 => (x"31",x"20",x"65",x"6c"),
  3963 => (x"2c",x"32",x"50",x"3b"),
  3964 => (x"74",x"73",x"79",x"53"),
  3965 => (x"50",x"3b",x"6d",x"65"),
  3966 => (x"4f",x"4e",x"4f",x"32"),
  3967 => (x"69",x"68",x"43",x"2c"),
  3968 => (x"74",x"65",x"73",x"70"),
  3969 => (x"2c",x"54",x"53",x"2c"),
  3970 => (x"2c",x"45",x"54",x"53"),
  3971 => (x"61",x"67",x"65",x"4d"),
  3972 => (x"2c",x"45",x"54",x"53"),
  3973 => (x"72",x"45",x"54",x"53"),
  3974 => (x"73",x"64",x"69",x"6f"),
  3975 => (x"4f",x"32",x"50",x"3b"),
  3976 => (x"54",x"53",x"2c",x"4a"),
  3977 => (x"69",x"6c",x"42",x"20"),
  3978 => (x"72",x"65",x"74",x"74"),
  3979 => (x"66",x"66",x"4f",x"2c"),
  3980 => (x"3b",x"6e",x"4f",x"2c"),
  3981 => (x"31",x"4f",x"32",x"50"),
  3982 => (x"41",x"52",x"2c",x"33"),
  3983 => (x"6e",x"28",x"20",x"4d"),
  3984 => (x"20",x"64",x"65",x"65"),
  3985 => (x"64",x"72",x"61",x"48"),
  3986 => (x"73",x"65",x"52",x"20"),
  3987 => (x"2c",x"29",x"74",x"65"),
  3988 => (x"4b",x"32",x"31",x"35"),
  3989 => (x"42",x"4d",x"31",x"2c"),
  3990 => (x"42",x"4d",x"32",x"2c"),
  3991 => (x"42",x"4d",x"34",x"2c"),
  3992 => (x"42",x"4d",x"38",x"2c"),
  3993 => (x"4d",x"34",x"31",x"2c"),
  3994 => (x"32",x"50",x"3b",x"42"),
  3995 => (x"4d",x"49",x"2c",x"46"),
  3996 => (x"4d",x"4f",x"52",x"47"),
  3997 => (x"61",x"6f",x"4c",x"2c"),
  3998 => (x"4f",x"52",x"20",x"64"),
  3999 => (x"32",x"50",x"3b",x"4d"),
  4000 => (x"49",x"42",x"2c",x"46"),
  4001 => (x"43",x"54",x"53",x"4e"),
  4002 => (x"61",x"6f",x"4c",x"2c"),
  4003 => (x"61",x"43",x"20",x"64"),
  4004 => (x"69",x"72",x"74",x"72"),
  4005 => (x"3b",x"65",x"67",x"64"),
  4006 => (x"53",x"2c",x"33",x"50"),
  4007 => (x"64",x"6e",x"75",x"6f"),
  4008 => (x"56",x"20",x"26",x"20"),
  4009 => (x"6f",x"65",x"64",x"69"),
  4010 => (x"4f",x"33",x"50",x"3b"),
  4011 => (x"69",x"56",x"2c",x"38"),
  4012 => (x"20",x"6f",x"65",x"64"),
  4013 => (x"65",x"64",x"6f",x"6d"),
  4014 => (x"6e",x"6f",x"4d",x"2c"),
  4015 => (x"6f",x"43",x"2c",x"6f"),
  4016 => (x"72",x"75",x"6f",x"6c"),
  4017 => (x"4f",x"33",x"50",x"3b"),
  4018 => (x"69",x"56",x"2c",x"53"),
  4019 => (x"67",x"6e",x"69",x"6b"),
  4020 => (x"31",x"4d",x"53",x"2f"),
  4021 => (x"4f",x"2c",x"34",x"39"),
  4022 => (x"4f",x"2c",x"66",x"66"),
  4023 => (x"33",x"50",x"3b",x"6e"),
  4024 => (x"2c",x"4c",x"4b",x"4f"),
  4025 => (x"6e",x"61",x"63",x"53"),
  4026 => (x"65",x"6e",x"69",x"6c"),
  4027 => (x"66",x"4f",x"2c",x"73"),
  4028 => (x"35",x"32",x"2c",x"66"),
  4029 => (x"30",x"35",x"2c",x"25"),
  4030 => (x"35",x"37",x"2c",x"25"),
  4031 => (x"33",x"50",x"3b",x"25"),
  4032 => (x"43",x"2c",x"54",x"4f"),
  4033 => (x"6f",x"70",x"6d",x"6f"),
  4034 => (x"65",x"74",x"69",x"73"),
  4035 => (x"65",x"6c",x"62",x"20"),
  4036 => (x"4f",x"2c",x"64",x"6e"),
  4037 => (x"4f",x"2c",x"66",x"66"),
  4038 => (x"33",x"50",x"3b",x"6e"),
  4039 => (x"53",x"2c",x"4d",x"4f"),
  4040 => (x"65",x"72",x"65",x"74"),
  4041 => (x"6f",x"73",x"20",x"6f"),
  4042 => (x"2c",x"64",x"6e",x"75"),
  4043 => (x"2c",x"66",x"66",x"4f"),
  4044 => (x"50",x"3b",x"6e",x"4f"),
  4045 => (x"2c",x"55",x"4f",x"33"),
  4046 => (x"69",x"65",x"74",x"53"),
  4047 => (x"72",x"65",x"62",x"6e"),
  4048 => (x"6f",x"64",x"20",x"67"),
  4049 => (x"65",x"6c",x"67",x"6e"),
  4050 => (x"66",x"66",x"4f",x"2c"),
  4051 => (x"3b",x"6e",x"4f",x"2c"),
  4052 => (x"43",x"2c",x"43",x"53"),
  4053 => (x"4c",x"2c",x"47",x"46"),
  4054 => (x"20",x"64",x"61",x"6f"),
  4055 => (x"66",x"6e",x"6f",x"63"),
  4056 => (x"53",x"3b",x"67",x"69"),
  4057 => (x"46",x"43",x"2c",x"44"),
  4058 => (x"61",x"53",x"2c",x"47"),
  4059 => (x"63",x"20",x"65",x"76"),
  4060 => (x"69",x"66",x"6e",x"6f"),
  4061 => (x"30",x"54",x"3b",x"67"),
  4062 => (x"73",x"65",x"52",x"2c"),
  4063 => (x"28",x"20",x"74",x"65"),
  4064 => (x"64",x"6c",x"6f",x"48"),
  4065 => (x"72",x"6f",x"66",x"20"),
  4066 => (x"72",x"61",x"68",x"20"),
  4067 => (x"65",x"72",x"20",x"64"),
  4068 => (x"29",x"74",x"65",x"73"),
  4069 => (x"76",x"2c",x"56",x"3b"),
  4070 => (x"30",x"34",x"2e",x"33"),
  4071 => (x"00",x"00",x"00",x"2e"),
  4072 => (x"20",x"53",x"4f",x"54"),
  4073 => (x"20",x"20",x"20",x"20"),
  4074 => (x"00",x"47",x"4d",x"49"),
  4075 => (x"54",x"53",x"49",x"4d"),
  4076 => (x"20",x"59",x"52",x"45"),
  4077 => (x"00",x"47",x"46",x"43"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

