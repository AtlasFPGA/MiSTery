library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0d9c487",
    12 => x"86c0c84e",
    13 => x"49c0d9c4",
    14 => x"48f8fec3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087fcf1",
    19 => x"fc1e87fd",
    20 => x"ff4a7186",
    21 => x"486949c0",
    22 => x"7098c0c4",
    23 => x"0298487e",
    24 => x"797287f4",
    25 => x"268efc48",
    26 => x"1e721e4f",
    27 => x"48121e73",
    28 => x"87ca0211",
    29 => x"98dfc34b",
    30 => x"0288739b",
    31 => x"4b2687f0",
    32 => x"4f264a26",
    33 => x"721e731e",
    34 => x"048bc11e",
    35 => x"481287ca",
    36 => x"87c40211",
    37 => x"87f10288",
    38 => x"4b264a26",
    39 => x"741e4f26",
    40 => x"721e731e",
    41 => x"048bc11e",
    42 => x"481287d0",
    43 => x"87ca0211",
    44 => x"98dfc34c",
    45 => x"0288749c",
    46 => x"4a2687eb",
    47 => x"4c264b26",
    48 => x"731e4f26",
    49 => x"a9738148",
    50 => x"1287c502",
    51 => x"87f60553",
    52 => x"731e4f26",
    53 => x"a9738148",
    54 => x"f9537205",
    55 => x"1e4f2687",
    56 => x"9a721e73",
    57 => x"87e7c002",
    58 => x"4bc148c0",
    59 => x"d106a972",
    60 => x"06827287",
    61 => x"837387c9",
    62 => x"f401a972",
    63 => x"c187c387",
    64 => x"a9723ab2",
    65 => x"80738903",
    66 => x"2b2ac107",
    67 => x"2687f305",
    68 => x"1e4f264b",
    69 => x"4dc41e75",
    70 => x"04a1b771",
    71 => x"81c1b9ff",
    72 => x"7207bdc3",
    73 => x"ff04a2b7",
    74 => x"c182c1ba",
    75 => x"eefe07bd",
    76 => x"042dc187",
    77 => x"80c1b8ff",
    78 => x"ff042d07",
    79 => x"0781c1b9",
    80 => x"4f264d26",
    81 => x"711e731e",
    82 => x"4b66c84a",
    83 => x"718bc149",
    84 => x"87cf0299",
    85 => x"d4ff4812",
    86 => x"49737808",
    87 => x"99718bc1",
    88 => x"2687f105",
    89 => x"0e4f264b",
    90 => x"0e5c5b5e",
    91 => x"d4ff4a71",
    92 => x"4b66cc4c",
    93 => x"718bc149",
    94 => x"87ce0299",
    95 => x"6c7cffc3",
    96 => x"c1497352",
    97 => x"0599718b",
    98 => x"4c2687f2",
    99 => x"4f264b26",
   100 => x"ff1e731e",
   101 => x"ffc34bd4",
   102 => x"c34a6b7b",
   103 => x"496b7bff",
   104 => x"b17232c8",
   105 => x"6b7bffc3",
   106 => x"7131c84a",
   107 => x"7bffc3b2",
   108 => x"32c8496b",
   109 => x"4871b172",
   110 => x"4f264b26",
   111 => x"5c5b5e0e",
   112 => x"4d710e5d",
   113 => x"754cd4ff",
   114 => x"98ffc348",
   115 => x"fec37c70",
   116 => x"c805bff8",
   117 => x"4866d087",
   118 => x"a6d430c9",
   119 => x"4966d058",
   120 => x"487129d8",
   121 => x"7098ffc3",
   122 => x"4966d07c",
   123 => x"487129d0",
   124 => x"7098ffc3",
   125 => x"4966d07c",
   126 => x"487129c8",
   127 => x"7098ffc3",
   128 => x"4866d07c",
   129 => x"7098ffc3",
   130 => x"d049757c",
   131 => x"c3487129",
   132 => x"7c7098ff",
   133 => x"f0c94b6c",
   134 => x"ffc34aff",
   135 => x"87cf05ab",
   136 => x"6c7c7149",
   137 => x"028ac14b",
   138 => x"ab7187c5",
   139 => x"7387f202",
   140 => x"264d2648",
   141 => x"264b264c",
   142 => x"49c01e4f",
   143 => x"c348d4ff",
   144 => x"81c178ff",
   145 => x"a9b7c8c3",
   146 => x"2687f104",
   147 => x"5b5e0e4f",
   148 => x"c00e5d5c",
   149 => x"f7c1f0ff",
   150 => x"c0c0c14d",
   151 => x"4bc0c0c0",
   152 => x"c487d6ff",
   153 => x"c04cdff8",
   154 => x"fd49751e",
   155 => x"86c487ce",
   156 => x"c005a8c1",
   157 => x"d4ff87e5",
   158 => x"78ffc348",
   159 => x"e1c01e73",
   160 => x"49e9c1f0",
   161 => x"c487f5fc",
   162 => x"05987086",
   163 => x"d4ff87ca",
   164 => x"78ffc348",
   165 => x"87cb48c1",
   166 => x"c187defe",
   167 => x"c6ff058c",
   168 => x"2648c087",
   169 => x"264c264d",
   170 => x"0e4f264b",
   171 => x"0e5c5b5e",
   172 => x"c1f0ffc0",
   173 => x"d4ff4cc1",
   174 => x"78ffc348",
   175 => x"1ec04bd3",
   176 => x"f7fb4974",
   177 => x"7086c487",
   178 => x"87ca0598",
   179 => x"c348d4ff",
   180 => x"48c178ff",
   181 => x"e0fd87ca",
   182 => x"058bc187",
   183 => x"48c087e0",
   184 => x"4b264c26",
   185 => x"5e0e4f26",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"c4fd4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"fbfa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087e0fe",
   195 => x"87e2c148",
   196 => x"7087fdf9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fe87c802",
   200 => x"48c087c9",
   201 => x"7587cbc1",
   202 => x"4cf1c07b",
   203 => x"7087defc",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87fcf949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"d548c187",
   215 => x"d148c087",
   216 => x"05acc287",
   217 => x"48c087c4",
   218 => x"8cc187c8",
   219 => x"87fcfe05",
   220 => x"4d2648c0",
   221 => x"4b264c26",
   222 => x"5e0e4f26",
   223 => x"0e5d5c5b",
   224 => x"c04dd0ff",
   225 => x"c0c1d0e5",
   226 => x"f8fec34c",
   227 => x"c778c148",
   228 => x"fa7dc24b",
   229 => x"7dc387e3",
   230 => x"49741ec0",
   231 => x"c487ddf8",
   232 => x"05a8c186",
   233 => x"c24b87c1",
   234 => x"87c505ab",
   235 => x"f6c048c0",
   236 => x"058bc187",
   237 => x"fc87daff",
   238 => x"fec387ec",
   239 => x"987058fc",
   240 => x"c187cd05",
   241 => x"f0ffc01e",
   242 => x"f749d0c1",
   243 => x"86c487ee",
   244 => x"c348d4ff",
   245 => x"e8c478ff",
   246 => x"c0ffc387",
   247 => x"ff7dc258",
   248 => x"ffc348d4",
   249 => x"2648c178",
   250 => x"264c264d",
   251 => x"0e4f264b",
   252 => x"5d5c5b5e",
   253 => x"c34d710e",
   254 => x"d4ff4cff",
   255 => x"ff7b744b",
   256 => x"c3c448d0",
   257 => x"757b7478",
   258 => x"f0ffc01e",
   259 => x"f649d8c1",
   260 => x"86c487ea",
   261 => x"c5029870",
   262 => x"c048c187",
   263 => x"7b7487ee",
   264 => x"c87bfec3",
   265 => x"66d41ec0",
   266 => x"87d8f449",
   267 => x"7b7486c4",
   268 => x"7b747b74",
   269 => x"4ae0dad8",
   270 => x"056b7b74",
   271 => x"8ac187c5",
   272 => x"7487f505",
   273 => x"48d0ff7b",
   274 => x"48c078c2",
   275 => x"4c264d26",
   276 => x"4f264b26",
   277 => x"5c5b5e0e",
   278 => x"86fc0e5d",
   279 => x"d4ff4b71",
   280 => x"c57ec04c",
   281 => x"4adfcdee",
   282 => x"6c7cffc3",
   283 => x"a8fec348",
   284 => x"87f8c005",
   285 => x"9b734d74",
   286 => x"d487cc02",
   287 => x"49731e66",
   288 => x"c487e4f3",
   289 => x"ff87d486",
   290 => x"d1c448d0",
   291 => x"4a66d478",
   292 => x"c17dffc3",
   293 => x"87f8058a",
   294 => x"c35aa6d8",
   295 => x"737c7cff",
   296 => x"87c5059b",
   297 => x"d048d0ff",
   298 => x"7e4ac178",
   299 => x"fe058ac1",
   300 => x"486e87f6",
   301 => x"4d268efc",
   302 => x"4b264c26",
   303 => x"731e4f26",
   304 => x"c04a711e",
   305 => x"48d4ff4b",
   306 => x"ff78ffc3",
   307 => x"c3c448d0",
   308 => x"48d4ff78",
   309 => x"7278ffc3",
   310 => x"f0ffc01e",
   311 => x"f349d1c1",
   312 => x"86c487da",
   313 => x"d2059870",
   314 => x"1ec0c887",
   315 => x"fd4966cc",
   316 => x"86c487e2",
   317 => x"d0ff4b70",
   318 => x"7378c248",
   319 => x"264b2648",
   320 => x"5b5e0e4f",
   321 => x"c00e5d5c",
   322 => x"f0ffc01e",
   323 => x"f249c9c1",
   324 => x"1ed287ea",
   325 => x"49c0ffc3",
   326 => x"c887f9fc",
   327 => x"c14cc086",
   328 => x"acb7d284",
   329 => x"c387f804",
   330 => x"bf97c0ff",
   331 => x"99c0c349",
   332 => x"05a9c0c1",
   333 => x"c387e7c0",
   334 => x"bf97c7ff",
   335 => x"c331d049",
   336 => x"bf97c8ff",
   337 => x"7232c84a",
   338 => x"c9ffc3b1",
   339 => x"b14abf97",
   340 => x"ffcf4c71",
   341 => x"c19cffff",
   342 => x"c134ca84",
   343 => x"ffc387e7",
   344 => x"49bf97c9",
   345 => x"99c631c1",
   346 => x"97caffc3",
   347 => x"b7c74abf",
   348 => x"c3b1722a",
   349 => x"bf97c5ff",
   350 => x"9dcf4d4a",
   351 => x"97c6ffc3",
   352 => x"9ac34abf",
   353 => x"ffc332ca",
   354 => x"4bbf97c7",
   355 => x"b27333c2",
   356 => x"97c8ffc3",
   357 => x"c0c34bbf",
   358 => x"2bb7c69b",
   359 => x"81c2b273",
   360 => x"307148c1",
   361 => x"48c14970",
   362 => x"4d703075",
   363 => x"84c14c72",
   364 => x"c0c89471",
   365 => x"cc06adb7",
   366 => x"b734c187",
   367 => x"b7c0c82d",
   368 => x"f4ff01ad",
   369 => x"26487487",
   370 => x"264c264d",
   371 => x"0e4f264b",
   372 => x"5d5c5b5e",
   373 => x"c486f80e",
   374 => x"c048e8c7",
   375 => x"e0ffc378",
   376 => x"fb49c01e",
   377 => x"86c487d8",
   378 => x"c5059870",
   379 => x"c948c087",
   380 => x"4dc087c0",
   381 => x"c2c17ec1",
   382 => x"c449bfd4",
   383 => x"714ad6c0",
   384 => x"ffe94bc8",
   385 => x"05987087",
   386 => x"7ec087c2",
   387 => x"bfd0c2c1",
   388 => x"f2c0c449",
   389 => x"4bc8714a",
   390 => x"7087e9e9",
   391 => x"87c20598",
   392 => x"026e7ec0",
   393 => x"c487fdc0",
   394 => x"4dbfe6c6",
   395 => x"9fdec7c4",
   396 => x"c5487ebf",
   397 => x"05a8ead6",
   398 => x"c6c487c7",
   399 => x"ce4dbfe6",
   400 => x"ca486e87",
   401 => x"02a8d5e9",
   402 => x"48c087c5",
   403 => x"c387e3c7",
   404 => x"751ee0ff",
   405 => x"87e6f949",
   406 => x"987086c4",
   407 => x"c087c505",
   408 => x"87cec748",
   409 => x"bfd0c2c1",
   410 => x"f2c0c449",
   411 => x"4bc8714a",
   412 => x"7087d1e8",
   413 => x"87c80598",
   414 => x"48e8c7c4",
   415 => x"87da78c1",
   416 => x"bfd4c2c1",
   417 => x"d6c0c449",
   418 => x"4bc8714a",
   419 => x"7087f5e7",
   420 => x"c5c00298",
   421 => x"c648c087",
   422 => x"c7c487d8",
   423 => x"49bf97de",
   424 => x"05a9d5c1",
   425 => x"c487cdc0",
   426 => x"bf97dfc7",
   427 => x"a9eac249",
   428 => x"87c5c002",
   429 => x"f9c548c0",
   430 => x"e0ffc387",
   431 => x"487ebf97",
   432 => x"02a8e9c3",
   433 => x"6e87cec0",
   434 => x"a8ebc348",
   435 => x"87c5c002",
   436 => x"ddc548c0",
   437 => x"ebffc387",
   438 => x"9949bf97",
   439 => x"87ccc005",
   440 => x"97ecffc3",
   441 => x"a9c249bf",
   442 => x"87c5c002",
   443 => x"c1c548c0",
   444 => x"edffc387",
   445 => x"c448bf97",
   446 => x"7058e4c7",
   447 => x"88c1484c",
   448 => x"58e8c7c4",
   449 => x"97eeffc3",
   450 => x"817549bf",
   451 => x"97efffc3",
   452 => x"32c84abf",
   453 => x"c47ea172",
   454 => x"6e48f8cb",
   455 => x"f0ffc378",
   456 => x"c848bf97",
   457 => x"c7c458a6",
   458 => x"c202bfe8",
   459 => x"c2c187cf",
   460 => x"c449bfd0",
   461 => x"714af2c0",
   462 => x"c7e54bc8",
   463 => x"02987087",
   464 => x"c087c5c0",
   465 => x"87eac348",
   466 => x"bfe0c7c4",
   467 => x"ccccc44c",
   468 => x"c5c0c45c",
   469 => x"c849bf97",
   470 => x"c4c0c431",
   471 => x"a14abf97",
   472 => x"c6c0c449",
   473 => x"d04abf97",
   474 => x"49a17232",
   475 => x"97c7c0c4",
   476 => x"32d84abf",
   477 => x"c449a172",
   478 => x"cbc49166",
   479 => x"c481bff8",
   480 => x"c459c0cc",
   481 => x"bf97cdc0",
   482 => x"c432c84a",
   483 => x"bf97ccc0",
   484 => x"c44aa24b",
   485 => x"bf97cec0",
   486 => x"7333d04b",
   487 => x"c0c44aa2",
   488 => x"4bbf97cf",
   489 => x"33d89bcf",
   490 => x"c44aa273",
   491 => x"c25ac4cc",
   492 => x"c492748a",
   493 => x"7248c4cc",
   494 => x"c1c178a1",
   495 => x"f2ffc387",
   496 => x"c849bf97",
   497 => x"f1ffc331",
   498 => x"a14abf97",
   499 => x"c731c549",
   500 => x"29c981ff",
   501 => x"59ccccc4",
   502 => x"97f7ffc3",
   503 => x"32c84abf",
   504 => x"97f6ffc3",
   505 => x"4aa24bbf",
   506 => x"6e9266c4",
   507 => x"c8ccc482",
   508 => x"c0ccc45a",
   509 => x"c478c048",
   510 => x"7248fccb",
   511 => x"ccc478a1",
   512 => x"ccc448cc",
   513 => x"c478bfc0",
   514 => x"c448d0cc",
   515 => x"78bfc4cc",
   516 => x"bfe8c7c4",
   517 => x"87c9c002",
   518 => x"30c44874",
   519 => x"c9c07e70",
   520 => x"c8ccc487",
   521 => x"30c448bf",
   522 => x"c7c47e70",
   523 => x"786e48ec",
   524 => x"8ef848c1",
   525 => x"4c264d26",
   526 => x"4f264b26",
   527 => x"5c5b5e0e",
   528 => x"4a710e5d",
   529 => x"bfe8c7c4",
   530 => x"7287cb02",
   531 => x"722bc74b",
   532 => x"9dffc14d",
   533 => x"4b7287c9",
   534 => x"4d722bc8",
   535 => x"c49dffc3",
   536 => x"83bff8cb",
   537 => x"bfccc2c1",
   538 => x"87d902ab",
   539 => x"5bd0c2c1",
   540 => x"1ee0ffc3",
   541 => x"c5f14973",
   542 => x"7086c487",
   543 => x"87c50598",
   544 => x"e6c048c0",
   545 => x"e8c7c487",
   546 => x"87d202bf",
   547 => x"91c44975",
   548 => x"81e0ffc3",
   549 => x"ffcf4c69",
   550 => x"9cffffff",
   551 => x"497587cb",
   552 => x"ffc391c2",
   553 => x"699f81e0",
   554 => x"2648744c",
   555 => x"264c264d",
   556 => x"0e4f264b",
   557 => x"5d5c5b5e",
   558 => x"cc86f00e",
   559 => x"66c859a6",
   560 => x"c087c505",
   561 => x"87c5c448",
   562 => x"c84866c8",
   563 => x"487e7080",
   564 => x"e0c078c0",
   565 => x"87c80266",
   566 => x"9766e0c0",
   567 => x"87c505bf",
   568 => x"e8c348c0",
   569 => x"c11ec087",
   570 => x"c4d14949",
   571 => x"7086c487",
   572 => x"c0029c4c",
   573 => x"c7c487fe",
   574 => x"e0c04af0",
   575 => x"ddff4966",
   576 => x"987087e7",
   577 => x"87ecc002",
   578 => x"e0c04a74",
   579 => x"4bcb4966",
   580 => x"87cadeff",
   581 => x"db029870",
   582 => x"741ec087",
   583 => x"87c4029c",
   584 => x"87c24dc0",
   585 => x"49754dc1",
   586 => x"c487c6d0",
   587 => x"9c4c7086",
   588 => x"87c2ff05",
   589 => x"c2029c74",
   590 => x"a4dc87d1",
   591 => x"69486e49",
   592 => x"49a4da78",
   593 => x"c44866c8",
   594 => x"58a6c880",
   595 => x"c448699f",
   596 => x"c4780866",
   597 => x"02bfe8c7",
   598 => x"a4d487d2",
   599 => x"49699f49",
   600 => x"99ffffc0",
   601 => x"30d04871",
   602 => x"87c558a6",
   603 => x"c048a6cc",
   604 => x"4966cc78",
   605 => x"bf66c448",
   606 => x"0866c480",
   607 => x"4866c878",
   608 => x"66c878c0",
   609 => x"c481cc49",
   610 => x"c879bf66",
   611 => x"81d04966",
   612 => x"c44d79c0",
   613 => x"66c84c66",
   614 => x"7582d44a",
   615 => x"7291c849",
   616 => x"41c049a1",
   617 => x"85c1796c",
   618 => x"04adb7c6",
   619 => x"6e87e7ff",
   620 => x"2ac94abf",
   621 => x"f0c04972",
   622 => x"e2dcff4a",
   623 => x"c84a7087",
   624 => x"c4c14966",
   625 => x"c1797281",
   626 => x"c087c248",
   627 => x"268ef048",
   628 => x"264c264d",
   629 => x"0e4f264b",
   630 => x"5d5c5b5e",
   631 => x"9c4c710e",
   632 => x"87cbc102",
   633 => x"6949a4c8",
   634 => x"87c3c102",
   635 => x"6c4a66d0",
   636 => x"48a6d049",
   637 => x"4d78a172",
   638 => x"e4c7c4b9",
   639 => x"baff4abf",
   640 => x"99719972",
   641 => x"87e4c002",
   642 => x"6b4ba4c4",
   643 => x"87ecf849",
   644 => x"c7c47b70",
   645 => x"6c49bfe0",
   646 => x"757c7181",
   647 => x"e4c7c4b9",
   648 => x"baff4abf",
   649 => x"99719972",
   650 => x"87dcff05",
   651 => x"267c66d0",
   652 => x"264c264d",
   653 => x"1e4f264b",
   654 => x"4b711e73",
   655 => x"87c7029b",
   656 => x"6949a3c8",
   657 => x"c087c505",
   658 => x"87f6c048",
   659 => x"bffccbc4",
   660 => x"4aa3c449",
   661 => x"8ac24a6a",
   662 => x"bfe0c7c4",
   663 => x"49a17292",
   664 => x"bfe4c7c4",
   665 => x"729a6b4a",
   666 => x"c2c149a1",
   667 => x"66c859d0",
   668 => x"c9e9711e",
   669 => x"7086c487",
   670 => x"87c40598",
   671 => x"87c248c0",
   672 => x"4b2648c1",
   673 => x"731e4f26",
   674 => x"9b4b711e",
   675 => x"c887c702",
   676 => x"056949a3",
   677 => x"48c087c5",
   678 => x"c487f6c0",
   679 => x"49bffccb",
   680 => x"6a4aa3c4",
   681 => x"c48ac24a",
   682 => x"92bfe0c7",
   683 => x"c449a172",
   684 => x"4abfe4c7",
   685 => x"a1729a6b",
   686 => x"d0c2c149",
   687 => x"1e66c859",
   688 => x"87ebe471",
   689 => x"987086c4",
   690 => x"c087c405",
   691 => x"c187c248",
   692 => x"264b2648",
   693 => x"5b5e0e4f",
   694 => x"f80e5d5c",
   695 => x"c47e7186",
   696 => x"78ff48a6",
   697 => x"ffffffc1",
   698 => x"c04dffff",
   699 => x"d44a6e4b",
   700 => x"c8497382",
   701 => x"49a17291",
   702 => x"694c66d8",
   703 => x"acb7c08c",
   704 => x"7587cb04",
   705 => x"c503acb7",
   706 => x"5ba6c887",
   707 => x"83c14d74",
   708 => x"04abb7c6",
   709 => x"c487d6ff",
   710 => x"8ef84866",
   711 => x"4c264d26",
   712 => x"4f264b26",
   713 => x"5c5b5e0e",
   714 => x"86f00e5d",
   715 => x"a6c47e71",
   716 => x"ffffc148",
   717 => x"78ffffff",
   718 => x"78ff80c4",
   719 => x"4cc04dc0",
   720 => x"83d44b6e",
   721 => x"92c84a74",
   722 => x"754aa273",
   723 => x"7391c849",
   724 => x"486a49a1",
   725 => x"a6d08869",
   726 => x"02ad7458",
   727 => x"66c487cf",
   728 => x"87c903a8",
   729 => x"c45ca6cc",
   730 => x"66cc48a6",
   731 => x"c684c178",
   732 => x"ff04acb7",
   733 => x"85c187ca",
   734 => x"04adb7c6",
   735 => x"c887fffe",
   736 => x"8ef04866",
   737 => x"4c264d26",
   738 => x"4f264b26",
   739 => x"5c5b5e0e",
   740 => x"86ec0e5d",
   741 => x"e4c04b71",
   742 => x"28c94866",
   743 => x"c458a6c8",
   744 => x"4abfe4c7",
   745 => x"4872baff",
   746 => x"cc9866c4",
   747 => x"9b7358a6",
   748 => x"87c1c302",
   749 => x"6949a3c8",
   750 => x"87f9c202",
   751 => x"986b4872",
   752 => x"c458a6d4",
   753 => x"7e6c4ca3",
   754 => x"d04866c8",
   755 => x"c605a866",
   756 => x"7b66c487",
   757 => x"c887ccc2",
   758 => x"49731e66",
   759 => x"c487f6fb",
   760 => x"c04d7086",
   761 => x"d004adb7",
   762 => x"4aa3d487",
   763 => x"91c84975",
   764 => x"2149a172",
   765 => x"c77c697b",
   766 => x"cc7bc087",
   767 => x"7c6949a3",
   768 => x"6b4866c4",
   769 => x"58a6c888",
   770 => x"731e66d0",
   771 => x"87c5fb49",
   772 => x"4d7086c4",
   773 => x"49a3c4c1",
   774 => x"6948a6c8",
   775 => x"4866d078",
   776 => x"06a866c8",
   777 => x"c087f2c0",
   778 => x"c004adb7",
   779 => x"a6cc87eb",
   780 => x"78a3d448",
   781 => x"91c84975",
   782 => x"d08166cc",
   783 => x"88694866",
   784 => x"66c84970",
   785 => x"87d106a9",
   786 => x"d7fb4973",
   787 => x"c8497087",
   788 => x"8166cc91",
   789 => x"6e4166d0",
   790 => x"1e66c479",
   791 => x"f6f54973",
   792 => x"c386c487",
   793 => x"731ee0ff",
   794 => x"87cbf749",
   795 => x"a3d086c4",
   796 => x"66e4c049",
   797 => x"268eec79",
   798 => x"264c264d",
   799 => x"1e4f264b",
   800 => x"4b711e73",
   801 => x"e4c0029b",
   802 => x"d0ccc487",
   803 => x"c24a735b",
   804 => x"e0c7c48a",
   805 => x"c49249bf",
   806 => x"48bffccb",
   807 => x"ccc48072",
   808 => x"487158d4",
   809 => x"c7c430c4",
   810 => x"edc058f0",
   811 => x"ccccc487",
   812 => x"c0ccc448",
   813 => x"ccc478bf",
   814 => x"ccc448d0",
   815 => x"c478bfc4",
   816 => x"02bfe8c7",
   817 => x"c7c487c9",
   818 => x"c449bfe0",
   819 => x"c487c731",
   820 => x"49bfc8cc",
   821 => x"c7c431c4",
   822 => x"4b2659f0",
   823 => x"c41e4f26",
   824 => x"49bfcccc",
   825 => x"bfc0ccc4",
   826 => x"87c405a9",
   827 => x"87c24ac0",
   828 => x"48724a71",
   829 => x"5e0e4f26",
   830 => x"710e5c5b",
   831 => x"724bc04a",
   832 => x"e1c0029a",
   833 => x"49a2da87",
   834 => x"c44b699f",
   835 => x"02bfe8c7",
   836 => x"a2d487cf",
   837 => x"49699f49",
   838 => x"ffffc04c",
   839 => x"c234d09c",
   840 => x"744cc087",
   841 => x"4973b349",
   842 => x"2687d4fd",
   843 => x"264b264c",
   844 => x"5b5e0e4f",
   845 => x"f00e5d5c",
   846 => x"59a6c886",
   847 => x"ffffffcf",
   848 => x"7ec04cf8",
   849 => x"d80266c4",
   850 => x"dcffc387",
   851 => x"c378c048",
   852 => x"c448d4ff",
   853 => x"78bfd0cc",
   854 => x"48d8ffc3",
   855 => x"bfccccc4",
   856 => x"fdc7c478",
   857 => x"c450c048",
   858 => x"49bfecc7",
   859 => x"bfdcffc3",
   860 => x"03aa714a",
   861 => x"7287ccc4",
   862 => x"0599cf49",
   863 => x"c187eac0",
   864 => x"c348ccc2",
   865 => x"78bfd4ff",
   866 => x"1ee0ffc3",
   867 => x"bfd4ffc3",
   868 => x"d4ffc349",
   869 => x"78a1c148",
   870 => x"e1dcff71",
   871 => x"c086c487",
   872 => x"c348e8fc",
   873 => x"cc78e0ff",
   874 => x"e8fcc087",
   875 => x"e0c048bf",
   876 => x"ecfcc080",
   877 => x"dcffc358",
   878 => x"80c148bf",
   879 => x"58e0ffc3",
   880 => x"000f2827",
   881 => x"bf97bf00",
   882 => x"c2029d4d",
   883 => x"e5c387e5",
   884 => x"dec202ad",
   885 => x"e8fcc087",
   886 => x"a3cb4bbf",
   887 => x"cf4c1149",
   888 => x"d2c105ac",
   889 => x"df497587",
   890 => x"cd89c199",
   891 => x"f0c7c491",
   892 => x"4aa3c181",
   893 => x"a3c35112",
   894 => x"c551124a",
   895 => x"51124aa3",
   896 => x"124aa3c7",
   897 => x"4aa3c951",
   898 => x"a3ce5112",
   899 => x"d051124a",
   900 => x"51124aa3",
   901 => x"124aa3d2",
   902 => x"4aa3d451",
   903 => x"a3d65112",
   904 => x"d851124a",
   905 => x"51124aa3",
   906 => x"124aa3dc",
   907 => x"4aa3de51",
   908 => x"7ec15112",
   909 => x"7487fcc0",
   910 => x"0599c849",
   911 => x"7487edc0",
   912 => x"0599d049",
   913 => x"e0c087d3",
   914 => x"ccc00266",
   915 => x"c0497387",
   916 => x"700f66e0",
   917 => x"d3c00298",
   918 => x"c0056e87",
   919 => x"c7c487c6",
   920 => x"50c048f0",
   921 => x"bfe8fcc0",
   922 => x"87ebc248",
   923 => x"48fdc7c4",
   924 => x"c47e50c0",
   925 => x"49bfecc7",
   926 => x"bfdcffc3",
   927 => x"04aa714a",
   928 => x"cf87f4fb",
   929 => x"f8ffffff",
   930 => x"d0ccc44c",
   931 => x"c8c005bf",
   932 => x"e8c7c487",
   933 => x"fcc102bf",
   934 => x"d8ffc387",
   935 => x"dbe649bf",
   936 => x"dcffc387",
   937 => x"48a6c458",
   938 => x"bfd8ffc3",
   939 => x"e8c7c478",
   940 => x"dbc002bf",
   941 => x"4966c487",
   942 => x"a9749974",
   943 => x"87c8c002",
   944 => x"c048a6c8",
   945 => x"87e7c078",
   946 => x"c148a6c8",
   947 => x"87dfc078",
   948 => x"cf4966c4",
   949 => x"a999f8ff",
   950 => x"87c8c002",
   951 => x"c048a6cc",
   952 => x"87c5c078",
   953 => x"c148a6cc",
   954 => x"48a6c878",
   955 => x"c87866cc",
   956 => x"e0c00566",
   957 => x"4966c487",
   958 => x"c7c489c2",
   959 => x"914abfe0",
   960 => x"bffccbc4",
   961 => x"d4ffc34a",
   962 => x"78a17248",
   963 => x"48dcffc3",
   964 => x"d2f978c0",
   965 => x"cf48c087",
   966 => x"f8ffffff",
   967 => x"268ef04c",
   968 => x"264c264d",
   969 => x"004f264b",
   970 => x"00000000",
   971 => x"5c5b5e0e",
   972 => x"86fc0e5d",
   973 => x"496e7e71",
   974 => x"c087c4f5",
   975 => x"4949c11e",
   976 => x"c487eef7",
   977 => x"9a4a7086",
   978 => x"87c7c102",
   979 => x"9f49a2da",
   980 => x"c7c44b69",
   981 => x"cf02bfe8",
   982 => x"49a2d487",
   983 => x"4c49699f",
   984 => x"9cffffc0",
   985 => x"87c234d0",
   986 => x"49744cc0",
   987 => x"66d44ba3",
   988 => x"87c405ab",
   989 => x"87dd48c1",
   990 => x"9a721ec0",
   991 => x"c087c402",
   992 => x"c187c24d",
   993 => x"f649754d",
   994 => x"86c487e7",
   995 => x"059a4a70",
   996 => x"c087f9fe",
   997 => x"268efc48",
   998 => x"264c264d",
   999 => x"0e4f264b",
  1000 => x"5d5c5b5e",
  1001 => x"c886f40e",
  1002 => x"66c459a6",
  1003 => x"4887c902",
  1004 => x"bfc0ccc4",
  1005 => x"87c505a8",
  1006 => x"f9c248c1",
  1007 => x"4966c487",
  1008 => x"c7c489c2",
  1009 => x"914abfe0",
  1010 => x"bffccbc4",
  1011 => x"c349a14a",
  1012 => x"711ee0ff",
  1013 => x"87e6d3ff",
  1014 => x"987086c4",
  1015 => x"c087c505",
  1016 => x"87d2c248",
  1017 => x"4ce0ffc3",
  1018 => x"6c977ec0",
  1019 => x"58a6cc48",
  1020 => x"c1029870",
  1021 => x"c34887ee",
  1022 => x"c102a8e5",
  1023 => x"a4cb87e6",
  1024 => x"49699749",
  1025 => x"c10299d0",
  1026 => x"4a7487da",
  1027 => x"49c0c2c1",
  1028 => x"c1ff4bc8",
  1029 => x"987087ee",
  1030 => x"87c8c105",
  1031 => x"c47ea4da",
  1032 => x"02bfe8c7",
  1033 => x"a4d487cf",
  1034 => x"49699f49",
  1035 => x"ffffc04d",
  1036 => x"c235d09d",
  1037 => x"6e4dc087",
  1038 => x"c849bf9f",
  1039 => x"a57148a6",
  1040 => x"dafd4978",
  1041 => x"02987087",
  1042 => x"66c487d4",
  1043 => x"4966cc1e",
  1044 => x"c487d9fb",
  1045 => x"02987086",
  1046 => x"7ec187c4",
  1047 => x"7ec087c2",
  1048 => x"87d2486e",
  1049 => x"6e84e0c0",
  1050 => x"7080c148",
  1051 => x"a8d0487e",
  1052 => x"87f6fd04",
  1053 => x"8ef448c0",
  1054 => x"4c264d26",
  1055 => x"4f264b26",
  1056 => x"20202e2e",
  1057 => x"20202020",
  1058 => x"00202020",
  1059 => x"ffffffff",
  1060 => x"00001098",
  1061 => x"000010a4",
  1062 => x"33544146",
  1063 => x"20202032",
  1064 => x"00000000",
  1065 => x"31544146",
  1066 => x"20202036",
  1067 => x"d0ff1e00",
  1068 => x"78e0c048",
  1069 => x"c21e4f26",
  1070 => x"7087ddd2",
  1071 => x"c6029949",
  1072 => x"a9fbc087",
  1073 => x"7187f005",
  1074 => x"0e4f2648",
  1075 => x"0e5c5b5e",
  1076 => x"4cc04b71",
  1077 => x"87c0d2c2",
  1078 => x"02994970",
  1079 => x"c087fac0",
  1080 => x"c002a9ec",
  1081 => x"fbc087f3",
  1082 => x"ecc002a9",
  1083 => x"b766cc87",
  1084 => x"87c703ac",
  1085 => x"c20266d0",
  1086 => x"71537187",
  1087 => x"87c20299",
  1088 => x"d1c284c1",
  1089 => x"497087d2",
  1090 => x"87cd0299",
  1091 => x"02a9ecc0",
  1092 => x"fbc087c7",
  1093 => x"d4ff05a9",
  1094 => x"0266d087",
  1095 => x"97c087c3",
  1096 => x"a9ecc07b",
  1097 => x"7487c405",
  1098 => x"7487c54a",
  1099 => x"8a0ac04a",
  1100 => x"4c264872",
  1101 => x"4f264b26",
  1102 => x"dbd0c21e",
  1103 => x"c04a7087",
  1104 => x"c904aaf0",
  1105 => x"aaf9c087",
  1106 => x"c087c301",
  1107 => x"c1c18af0",
  1108 => x"87c904aa",
  1109 => x"01aadac1",
  1110 => x"f7c087c3",
  1111 => x"2648728a",
  1112 => x"5b5e0e4f",
  1113 => x"f80e5d5c",
  1114 => x"c04c7186",
  1115 => x"cad0c27e",
  1116 => x"c14bc087",
  1117 => x"bf97c4c8",
  1118 => x"04a9c049",
  1119 => x"f5fc87cf",
  1120 => x"c183c187",
  1121 => x"bf97c4c8",
  1122 => x"f106ab49",
  1123 => x"c4c8c187",
  1124 => x"d002bf97",
  1125 => x"ffcec287",
  1126 => x"99497087",
  1127 => x"c087c602",
  1128 => x"f005a9ec",
  1129 => x"c24bc087",
  1130 => x"7087edce",
  1131 => x"e7cec24d",
  1132 => x"58a6c887",
  1133 => x"87e0cec2",
  1134 => x"83c14a70",
  1135 => x"9749a4c8",
  1136 => x"05ad4969",
  1137 => x"a4c987da",
  1138 => x"49699749",
  1139 => x"05a966c4",
  1140 => x"a4ca87ce",
  1141 => x"49699749",
  1142 => x"87c405aa",
  1143 => x"87d07ec1",
  1144 => x"02adecc0",
  1145 => x"fbc087c6",
  1146 => x"87c405ad",
  1147 => x"7ec14bc0",
  1148 => x"f2fe026e",
  1149 => x"87f5fa87",
  1150 => x"8ef84873",
  1151 => x"4c264d26",
  1152 => x"4f264b26",
  1153 => x"5b5e0e00",
  1154 => x"f40e5d5c",
  1155 => x"ff7e7186",
  1156 => x"1e6e4bd4",
  1157 => x"49dcccc4",
  1158 => x"87d7daff",
  1159 => x"987086c4",
  1160 => x"87f7c402",
  1161 => x"c148a6c4",
  1162 => x"78bfe8f3",
  1163 => x"f0fc496e",
  1164 => x"58a6cc87",
  1165 => x"c5059870",
  1166 => x"48a6c887",
  1167 => x"d0ff78c1",
  1168 => x"c178c548",
  1169 => x"66c87bd5",
  1170 => x"c689c149",
  1171 => x"e0f3c131",
  1172 => x"484abf97",
  1173 => x"7b70b071",
  1174 => x"c448d0ff",
  1175 => x"d4ccc478",
  1176 => x"d049bf97",
  1177 => x"87d70299",
  1178 => x"d6c178c5",
  1179 => x"c34ac07b",
  1180 => x"82c17bff",
  1181 => x"04aae0c0",
  1182 => x"d0ff87f5",
  1183 => x"c378c448",
  1184 => x"d0ff7bff",
  1185 => x"c178c548",
  1186 => x"7bc17bd3",
  1187 => x"7e7378c4",
  1188 => x"c04866c4",
  1189 => x"c206a8b7",
  1190 => x"ccc487ee",
  1191 => x"c44cbfe4",
  1192 => x"88744866",
  1193 => x"7458a6c8",
  1194 => x"f7c1029c",
  1195 => x"e0ffc387",
  1196 => x"4bc0c84d",
  1197 => x"acb7c08c",
  1198 => x"c887c603",
  1199 => x"c04ba4c0",
  1200 => x"d4ccc44c",
  1201 => x"d049bf97",
  1202 => x"87d10299",
  1203 => x"ccc41ec0",
  1204 => x"ddff49dc",
  1205 => x"86c487e1",
  1206 => x"ebc04a70",
  1207 => x"e0ffc387",
  1208 => x"dcccc41e",
  1209 => x"ceddff49",
  1210 => x"7086c487",
  1211 => x"48d0ff4a",
  1212 => x"6e78c5c8",
  1213 => x"78d4c148",
  1214 => x"086e4815",
  1215 => x"058bc178",
  1216 => x"ff87f5ff",
  1217 => x"78c448d0",
  1218 => x"c5059a72",
  1219 => x"c148c087",
  1220 => x"1ec187cb",
  1221 => x"49dcccc4",
  1222 => x"87fbdaff",
  1223 => x"9c7486c4",
  1224 => x"87c9fe05",
  1225 => x"c04866c4",
  1226 => x"d106a8b7",
  1227 => x"dcccc487",
  1228 => x"d078c048",
  1229 => x"f478c080",
  1230 => x"e8ccc480",
  1231 => x"66c478bf",
  1232 => x"a8b7c048",
  1233 => x"87d2fd01",
  1234 => x"d0ff4b6e",
  1235 => x"c178c548",
  1236 => x"7bc07bd3",
  1237 => x"48c178c4",
  1238 => x"c087c2c0",
  1239 => x"268ef448",
  1240 => x"264c264d",
  1241 => x"0e4f264b",
  1242 => x"5d5c5b5e",
  1243 => x"7186fc0e",
  1244 => x"4c4bc04d",
  1245 => x"e8c004ad",
  1246 => x"e1c5c187",
  1247 => x"029c741e",
  1248 => x"4ac087c4",
  1249 => x"4ac187c2",
  1250 => x"e4e64972",
  1251 => x"7086c487",
  1252 => x"6e83c17e",
  1253 => x"7587c205",
  1254 => x"7584c14b",
  1255 => x"d8ff06ab",
  1256 => x"fc486e87",
  1257 => x"264d268e",
  1258 => x"264b264c",
  1259 => x"5b5e0e4f",
  1260 => x"fc0e5d5c",
  1261 => x"494c7186",
  1262 => x"cdc491de",
  1263 => x"85714df8",
  1264 => x"c1026d97",
  1265 => x"cdc487dd",
  1266 => x"7449bfe4",
  1267 => x"d6fe7181",
  1268 => x"487e7087",
  1269 => x"f3c00298",
  1270 => x"eccdc487",
  1271 => x"cb4a704b",
  1272 => x"ddf3fe49",
  1273 => x"cc4b7487",
  1274 => x"fcf3c193",
  1275 => x"c183c483",
  1276 => x"747bf0d0",
  1277 => x"e7c6c149",
  1278 => x"c17b7587",
  1279 => x"bf97e4f3",
  1280 => x"cdc41e49",
  1281 => x"d5c249ec",
  1282 => x"86c487d6",
  1283 => x"c6c14974",
  1284 => x"49c087ce",
  1285 => x"87e9c7c1",
  1286 => x"48d8ccc4",
  1287 => x"49c178c0",
  1288 => x"fc87c4de",
  1289 => x"264d268e",
  1290 => x"264b264c",
  1291 => x"0000004f",
  1292 => x"64616f4c",
  1293 => x"2e676e69",
  1294 => x"1e002e2e",
  1295 => x"4a711e73",
  1296 => x"e4cdc449",
  1297 => x"fc7181bf",
  1298 => x"4b7087dd",
  1299 => x"87c4029b",
  1300 => x"87e2e249",
  1301 => x"48e4cdc4",
  1302 => x"49c178c0",
  1303 => x"2687c8dd",
  1304 => x"1e4f264b",
  1305 => x"c6c149c0",
  1306 => x"4f2687d7",
  1307 => x"494a711e",
  1308 => x"f3c191cc",
  1309 => x"81c881fc",
  1310 => x"ccc44811",
  1311 => x"cdc458dc",
  1312 => x"78c048e4",
  1313 => x"dedc49c1",
  1314 => x"1e4f2687",
  1315 => x"d2029971",
  1316 => x"d8f5c187",
  1317 => x"f750c048",
  1318 => x"ecd1c180",
  1319 => x"f4f3c140",
  1320 => x"c187ce78",
  1321 => x"c148d4f5",
  1322 => x"fc78ecf3",
  1323 => x"e3d1c180",
  1324 => x"0e4f2678",
  1325 => x"5d5c5b5e",
  1326 => x"c386f40e",
  1327 => x"c04de0ff",
  1328 => x"48a6c84c",
  1329 => x"7e7578c0",
  1330 => x"bfe4cdc4",
  1331 => x"06a8c048",
  1332 => x"c887c0c1",
  1333 => x"7e755ca6",
  1334 => x"48e0ffc3",
  1335 => x"f2c00298",
  1336 => x"4d66c487",
  1337 => x"1ee1c5c1",
  1338 => x"c40266cc",
  1339 => x"c24cc087",
  1340 => x"744cc187",
  1341 => x"87f9e049",
  1342 => x"7e7086c4",
  1343 => x"66c885c1",
  1344 => x"cc80c148",
  1345 => x"cdc458a6",
  1346 => x"03adbfe4",
  1347 => x"056e87c5",
  1348 => x"6e87d1ff",
  1349 => x"754cc04d",
  1350 => x"ddc3029d",
  1351 => x"e1c5c187",
  1352 => x"0266cc1e",
  1353 => x"a6c887c7",
  1354 => x"c578c048",
  1355 => x"48a6c887",
  1356 => x"66c878c1",
  1357 => x"f8dfff49",
  1358 => x"7086c487",
  1359 => x"0298487e",
  1360 => x"4987e4c2",
  1361 => x"699781cb",
  1362 => x"0299d049",
  1363 => x"7487d4c1",
  1364 => x"c191cc49",
  1365 => x"c181fcf3",
  1366 => x"c879fbd0",
  1367 => x"51ffc381",
  1368 => x"91de4974",
  1369 => x"4df8cdc4",
  1370 => x"c1c28571",
  1371 => x"a5c17d97",
  1372 => x"51e0c049",
  1373 => x"97f0c7c4",
  1374 => x"87d202bf",
  1375 => x"a5c284c1",
  1376 => x"f0c7c44b",
  1377 => x"fe49db4a",
  1378 => x"c187f7ec",
  1379 => x"a5cd87d9",
  1380 => x"c151c049",
  1381 => x"4ba5c284",
  1382 => x"49cb4a6e",
  1383 => x"87e2ecfe",
  1384 => x"7487c4c1",
  1385 => x"c191cc49",
  1386 => x"c181fcf3",
  1387 => x"c479edce",
  1388 => x"bf97f0c7",
  1389 => x"7487d802",
  1390 => x"c191de49",
  1391 => x"f8cdc484",
  1392 => x"c483714b",
  1393 => x"dd4af0c7",
  1394 => x"f5ebfe49",
  1395 => x"7487d887",
  1396 => x"c493de4b",
  1397 => x"cb83f8cd",
  1398 => x"51c049a3",
  1399 => x"6e7384c1",
  1400 => x"fe49cb4a",
  1401 => x"c887dbeb",
  1402 => x"80c14866",
  1403 => x"c758a6cc",
  1404 => x"c5c003ac",
  1405 => x"fc056e87",
  1406 => x"487487e3",
  1407 => x"4d268ef4",
  1408 => x"4b264c26",
  1409 => x"731e4f26",
  1410 => x"494b711e",
  1411 => x"f3c191cc",
  1412 => x"a1c881fc",
  1413 => x"e0f3c14a",
  1414 => x"c9501248",
  1415 => x"c8c14aa1",
  1416 => x"501248c4",
  1417 => x"f3c181ca",
  1418 => x"501148e4",
  1419 => x"97e4f3c1",
  1420 => x"c01e49bf",
  1421 => x"e7ccc249",
  1422 => x"d8ccc487",
  1423 => x"c178de48",
  1424 => x"87e3d549",
  1425 => x"4b268efc",
  1426 => x"5e0e4f26",
  1427 => x"0e5d5c5b",
  1428 => x"4d7186f4",
  1429 => x"c191cc49",
  1430 => x"c881fcf3",
  1431 => x"a1ca4aa1",
  1432 => x"48a6c47e",
  1433 => x"bff4d1c4",
  1434 => x"bf976e78",
  1435 => x"4c66c44b",
  1436 => x"48122c73",
  1437 => x"7058a6cc",
  1438 => x"c984c19c",
  1439 => x"49699781",
  1440 => x"c204acb7",
  1441 => x"6e4cc087",
  1442 => x"c84abf97",
  1443 => x"31724966",
  1444 => x"66c4b9ff",
  1445 => x"72487499",
  1446 => x"484a7030",
  1447 => x"d1c4b071",
  1448 => x"f9c158f8",
  1449 => x"49c087f9",
  1450 => x"7587fcd3",
  1451 => x"effbc049",
  1452 => x"268ef487",
  1453 => x"264c264d",
  1454 => x"1e4f264b",
  1455 => x"4b711e73",
  1456 => x"024aa3c6",
  1457 => x"8ac187db",
  1458 => x"8a87d602",
  1459 => x"87dac102",
  1460 => x"fcc0028a",
  1461 => x"c0028a87",
  1462 => x"028a87e1",
  1463 => x"dbc187cb",
  1464 => x"f649c787",
  1465 => x"dec187c6",
  1466 => x"e4cdc487",
  1467 => x"cbc102bf",
  1468 => x"88c14887",
  1469 => x"58e8cdc4",
  1470 => x"c487c1c1",
  1471 => x"02bfe8cd",
  1472 => x"c487f9c0",
  1473 => x"48bfe4cd",
  1474 => x"cdc480c1",
  1475 => x"ebc058e8",
  1476 => x"e4cdc487",
  1477 => x"89c649bf",
  1478 => x"59e8cdc4",
  1479 => x"03a9b7c0",
  1480 => x"cdc487da",
  1481 => x"78c048e4",
  1482 => x"cdc487d2",
  1483 => x"cb02bfe8",
  1484 => x"e4cdc487",
  1485 => x"80c648bf",
  1486 => x"58e8cdc4",
  1487 => x"e6d149c0",
  1488 => x"c0497387",
  1489 => x"2687d9f9",
  1490 => x"0e4f264b",
  1491 => x"5d5c5b5e",
  1492 => x"86d4ff0e",
  1493 => x"c859a6dc",
  1494 => x"78c048a6",
  1495 => x"c0c180c4",
  1496 => x"80c47866",
  1497 => x"80c478c1",
  1498 => x"cdc478c1",
  1499 => x"78c148e8",
  1500 => x"bfd8ccc4",
  1501 => x"05a8de48",
  1502 => x"f6f487c9",
  1503 => x"58a6cc87",
  1504 => x"c187dfcf",
  1505 => x"e487f4f7",
  1506 => x"f7c187ec",
  1507 => x"4c7087ca",
  1508 => x"02acfbc0",
  1509 => x"d887f0c1",
  1510 => x"e2c10566",
  1511 => x"66fcc087",
  1512 => x"6a82c44a",
  1513 => x"d8eec17e",
  1514 => x"20496e48",
  1515 => x"10412041",
  1516 => x"66fcc051",
  1517 => x"c6d8c148",
  1518 => x"c7496a78",
  1519 => x"c0517481",
  1520 => x"c84966fc",
  1521 => x"c051c181",
  1522 => x"c94966fc",
  1523 => x"c051c081",
  1524 => x"ca4966fc",
  1525 => x"c151c081",
  1526 => x"6a1ed81e",
  1527 => x"e381c849",
  1528 => x"86c887e9",
  1529 => x"4866c0c1",
  1530 => x"c701a8c0",
  1531 => x"48a6c887",
  1532 => x"87ce78c1",
  1533 => x"4866c0c1",
  1534 => x"a6d088c1",
  1535 => x"e287c358",
  1536 => x"a6d087f4",
  1537 => x"7478c248",
  1538 => x"d1cd029c",
  1539 => x"4866c887",
  1540 => x"a866c4c1",
  1541 => x"87c6cd03",
  1542 => x"c048a6dc",
  1543 => x"f4c17e78",
  1544 => x"4c7087f6",
  1545 => x"05acd0c1",
  1546 => x"c487d9c2",
  1547 => x"786e48a6",
  1548 => x"7087c5e4",
  1549 => x"dff4c17e",
  1550 => x"c04c7087",
  1551 => x"c105acec",
  1552 => x"66c887ed",
  1553 => x"c091cc49",
  1554 => x"c48166fc",
  1555 => x"4d6a4aa1",
  1556 => x"6e4aa1c8",
  1557 => x"ecd1c152",
  1558 => x"fbf3c179",
  1559 => x"9c4c7087",
  1560 => x"c087d902",
  1561 => x"d302acfb",
  1562 => x"c1557487",
  1563 => x"7087e9f3",
  1564 => x"c7029c4c",
  1565 => x"acfbc087",
  1566 => x"87edff05",
  1567 => x"c255e0c0",
  1568 => x"97c055c1",
  1569 => x"4866d87d",
  1570 => x"05a866c4",
  1571 => x"66c887db",
  1572 => x"a866cc48",
  1573 => x"c887ca04",
  1574 => x"80c14866",
  1575 => x"c858a6cc",
  1576 => x"4866cc87",
  1577 => x"a6d088c1",
  1578 => x"ebf2c158",
  1579 => x"c14c7087",
  1580 => x"c805acd0",
  1581 => x"4866d487",
  1582 => x"a6d880c1",
  1583 => x"acd0c158",
  1584 => x"87e7fd02",
  1585 => x"66d8486e",
  1586 => x"e3c905a8",
  1587 => x"a6e0c087",
  1588 => x"7478c048",
  1589 => x"88fbc048",
  1590 => x"7058a6c8",
  1591 => x"e4c90298",
  1592 => x"88cb4887",
  1593 => x"7058a6c8",
  1594 => x"d1c10298",
  1595 => x"88c94887",
  1596 => x"7058a6c8",
  1597 => x"c1c40298",
  1598 => x"88c44887",
  1599 => x"7058a6c8",
  1600 => x"87cf0298",
  1601 => x"c888c148",
  1602 => x"987058a6",
  1603 => x"87eac302",
  1604 => x"dc87d4c8",
  1605 => x"f0c048a6",
  1606 => x"fbf0c178",
  1607 => x"c04c7087",
  1608 => x"c002acec",
  1609 => x"e0c087c4",
  1610 => x"ecc05ca6",
  1611 => x"cdc002ac",
  1612 => x"e3f0c187",
  1613 => x"c04c7087",
  1614 => x"ff05acec",
  1615 => x"ecc087f3",
  1616 => x"c4c002ac",
  1617 => x"cff0c187",
  1618 => x"ca1ec087",
  1619 => x"4966d01e",
  1620 => x"c4c191cc",
  1621 => x"80714866",
  1622 => x"c858a6cc",
  1623 => x"80c44866",
  1624 => x"cc58a6d0",
  1625 => x"ff49bf66",
  1626 => x"c187e0dd",
  1627 => x"d41ede1e",
  1628 => x"ff49bf66",
  1629 => x"d087d4dd",
  1630 => x"48497086",
  1631 => x"c08808c0",
  1632 => x"c058a6e8",
  1633 => x"eec006a8",
  1634 => x"66e4c087",
  1635 => x"03a8dd48",
  1636 => x"c487e4c0",
  1637 => x"c049bf66",
  1638 => x"c08166e4",
  1639 => x"e4c051e0",
  1640 => x"81c14966",
  1641 => x"81bf66c4",
  1642 => x"c051c1c2",
  1643 => x"c24966e4",
  1644 => x"bf66c481",
  1645 => x"6e51c081",
  1646 => x"c6d8c148",
  1647 => x"c8496e78",
  1648 => x"5166d081",
  1649 => x"81c9496e",
  1650 => x"6e5166d4",
  1651 => x"dc81ca49",
  1652 => x"66d05166",
  1653 => x"d480c148",
  1654 => x"66c858a6",
  1655 => x"a866cc48",
  1656 => x"87cbc004",
  1657 => x"c14866c8",
  1658 => x"58a6cc80",
  1659 => x"cc87d6c5",
  1660 => x"88c14866",
  1661 => x"c558a6d0",
  1662 => x"dcff87cb",
  1663 => x"e8c087fa",
  1664 => x"dcff58a6",
  1665 => x"e0c087f2",
  1666 => x"ecc058a6",
  1667 => x"cac005a8",
  1668 => x"48a6dc87",
  1669 => x"7866e4c0",
  1670 => x"c187c4c0",
  1671 => x"c887f9ec",
  1672 => x"91cc4966",
  1673 => x"4866fcc0",
  1674 => x"a6c88071",
  1675 => x"4a66c458",
  1676 => x"66c482c8",
  1677 => x"c081ca49",
  1678 => x"dc5166e4",
  1679 => x"81c14966",
  1680 => x"8966e4c0",
  1681 => x"307148c1",
  1682 => x"89c14970",
  1683 => x"c47a9771",
  1684 => x"49bff4d1",
  1685 => x"2966e4c0",
  1686 => x"484a6a97",
  1687 => x"ecc09871",
  1688 => x"66c458a6",
  1689 => x"6981c449",
  1690 => x"4866d84d",
  1691 => x"c002a86e",
  1692 => x"7ec087c5",
  1693 => x"c187c2c0",
  1694 => x"c01e6e7e",
  1695 => x"49751ee0",
  1696 => x"87c7d9ff",
  1697 => x"4c7086c8",
  1698 => x"06acb7c0",
  1699 => x"7487d0c1",
  1700 => x"49e0c085",
  1701 => x"4b758974",
  1702 => x"4ae4eec1",
  1703 => x"e1d8fe71",
  1704 => x"7585c287",
  1705 => x"66e0c07e",
  1706 => x"c080c148",
  1707 => x"c058a6e4",
  1708 => x"c14966e8",
  1709 => x"02a97081",
  1710 => x"c087c5c0",
  1711 => x"87c2c04d",
  1712 => x"1e754dc1",
  1713 => x"c049a4c2",
  1714 => x"887148e0",
  1715 => x"c81e4970",
  1716 => x"d7ff4966",
  1717 => x"86c887f5",
  1718 => x"01a8b7c0",
  1719 => x"c087c6ff",
  1720 => x"c00266e0",
  1721 => x"66c487d3",
  1722 => x"c081c949",
  1723 => x"c45166e0",
  1724 => x"d9c14866",
  1725 => x"cec078ca",
  1726 => x"4966c487",
  1727 => x"51c281c9",
  1728 => x"c34866c4",
  1729 => x"c878d8dd",
  1730 => x"66cc4866",
  1731 => x"cbc004a8",
  1732 => x"4866c887",
  1733 => x"a6cc80c1",
  1734 => x"87e9c058",
  1735 => x"c14866cc",
  1736 => x"58a6d088",
  1737 => x"ff87dec0",
  1738 => x"7087cbd6",
  1739 => x"87d5c04c",
  1740 => x"05acc6c1",
  1741 => x"d087c8c0",
  1742 => x"80c14866",
  1743 => x"ff58a6d4",
  1744 => x"7087f3d5",
  1745 => x"4866d44c",
  1746 => x"a6d880c1",
  1747 => x"029c7458",
  1748 => x"c887cbc0",
  1749 => x"c4c14866",
  1750 => x"f204a866",
  1751 => x"d5ff87fa",
  1752 => x"66c887cb",
  1753 => x"03a8c748",
  1754 => x"c887e1c0",
  1755 => x"cdc44c66",
  1756 => x"78c048e8",
  1757 => x"91cc4974",
  1758 => x"8166fcc0",
  1759 => x"6a4aa1c4",
  1760 => x"7952c04a",
  1761 => x"acc784c1",
  1762 => x"87e2ff04",
  1763 => x"268ed4ff",
  1764 => x"264c264d",
  1765 => x"004f264b",
  1766 => x"64616f4c",
  1767 => x"202e2a20",
  1768 => x"00000000",
  1769 => x"1e00203a",
  1770 => x"4b711e73",
  1771 => x"87c6029b",
  1772 => x"48e4cdc4",
  1773 => x"1ec778c0",
  1774 => x"bfe4cdc4",
  1775 => x"fcf3c11e",
  1776 => x"d8ccc41e",
  1777 => x"c2ee49bf",
  1778 => x"c486cc87",
  1779 => x"49bfd8cc",
  1780 => x"7387f8e2",
  1781 => x"87c8029b",
  1782 => x"49fcf3c1",
  1783 => x"87cee8c0",
  1784 => x"4f264b26",
  1785 => x"fc1e731e",
  1786 => x"4bffc386",
  1787 => x"fc4ad4ff",
  1788 => x"98c148bf",
  1789 => x"98487e70",
  1790 => x"87fbc002",
  1791 => x"c148d0ff",
  1792 => x"d2c278c1",
  1793 => x"c37a737a",
  1794 => x"4849e1ff",
  1795 => x"506a80ff",
  1796 => x"516a7a73",
  1797 => x"80c17a73",
  1798 => x"7a73506a",
  1799 => x"7a73506a",
  1800 => x"7a73496a",
  1801 => x"7a73506a",
  1802 => x"ffc3506a",
  1803 => x"ff5997ea",
  1804 => x"c0c148d0",
  1805 => x"c387d778",
  1806 => x"4849e1ff",
  1807 => x"50c080ff",
  1808 => x"c080c151",
  1809 => x"c150d950",
  1810 => x"50e2c050",
  1811 => x"ffc350c3",
  1812 => x"50c048e7",
  1813 => x"8efc80f8",
  1814 => x"4f264b26",
  1815 => x"87d5cc1e",
  1816 => x"c2fd49c1",
  1817 => x"d1dcfe87",
  1818 => x"02987087",
  1819 => x"e5fe87cd",
  1820 => x"987087dd",
  1821 => x"c187c402",
  1822 => x"c087c24a",
  1823 => x"059a724a",
  1824 => x"1ec087ce",
  1825 => x"49f0f2c1",
  1826 => x"87edf2c0",
  1827 => x"87fe86c4",
  1828 => x"f2c11ec0",
  1829 => x"f2c049fc",
  1830 => x"1ec087df",
  1831 => x"87d1f9c1",
  1832 => x"f2c04970",
  1833 => x"d7c387d3",
  1834 => x"268ef887",
  1835 => x"0000004f",
  1836 => x"66204453",
  1837 => x"656c6961",
  1838 => x"00002e64",
  1839 => x"746f6f42",
  1840 => x"2e676e69",
  1841 => x"1e002e2e",
  1842 => x"48e4cdc4",
  1843 => x"ccc478c0",
  1844 => x"78c048d8",
  1845 => x"c187c5fe",
  1846 => x"c087f3fb",
  1847 => x"004f2648",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000001",
  1851 => x"78452080",
  1852 => x"00007469",
  1853 => x"61422080",
  1854 => x"00006b63",
  1855 => x"000013ad",
  1856 => x"00004378",
  1857 => x"00000000",
  1858 => x"000013ad",
  1859 => x"00004396",
  1860 => x"00000000",
  1861 => x"000013ad",
  1862 => x"000043b4",
  1863 => x"00000000",
  1864 => x"000013ad",
  1865 => x"000043d2",
  1866 => x"00000000",
  1867 => x"000013ad",
  1868 => x"000043f0",
  1869 => x"00000000",
  1870 => x"000013ad",
  1871 => x"0000440e",
  1872 => x"00000000",
  1873 => x"000013ad",
  1874 => x"0000442c",
  1875 => x"00000000",
  1876 => x"0000146c",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"000016bb",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"48f0fe1e",
  1883 => x"09cd78c0",
  1884 => x"4f260979",
  1885 => x"fe86fc1e",
  1886 => x"487ebff0",
  1887 => x"4f268efc",
  1888 => x"48f0fe1e",
  1889 => x"4f2678c1",
  1890 => x"48f0fe1e",
  1891 => x"4f2678c0",
  1892 => x"c04a711e",
  1893 => x"a2c17a97",
  1894 => x"ca51c049",
  1895 => x"51c049a2",
  1896 => x"c049a2cb",
  1897 => x"0e4f2651",
  1898 => x"0e5c5b5e",
  1899 => x"4c7186f0",
  1900 => x"9749a4ca",
  1901 => x"a4cb7e69",
  1902 => x"486b974b",
  1903 => x"c158a6c8",
  1904 => x"58a6cc80",
  1905 => x"a6d098c7",
  1906 => x"cc486e58",
  1907 => x"db05a866",
  1908 => x"7e699787",
  1909 => x"c8486b97",
  1910 => x"80c158a6",
  1911 => x"c758a6cc",
  1912 => x"58a6d098",
  1913 => x"66cc486e",
  1914 => x"87e502a8",
  1915 => x"cc87d9fe",
  1916 => x"6b974aa4",
  1917 => x"49a17249",
  1918 => x"975166dc",
  1919 => x"486e7e6b",
  1920 => x"a6c880c1",
  1921 => x"cc98c758",
  1922 => x"977058a6",
  1923 => x"87d1c27b",
  1924 => x"f087edfd",
  1925 => x"264c268e",
  1926 => x"0e4f264b",
  1927 => x"5d5c5b5e",
  1928 => x"7186f40e",
  1929 => x"7e6d974d",
  1930 => x"974ca5c1",
  1931 => x"a6c8486c",
  1932 => x"c4486e58",
  1933 => x"c505a866",
  1934 => x"c048ff87",
  1935 => x"c7fd87e6",
  1936 => x"49a5c287",
  1937 => x"714b6c97",
  1938 => x"6b974ba3",
  1939 => x"7e6c974b",
  1940 => x"80c1486e",
  1941 => x"c758a6c8",
  1942 => x"58a6cc98",
  1943 => x"fc7c9770",
  1944 => x"487387de",
  1945 => x"4d268ef4",
  1946 => x"4b264c26",
  1947 => x"5e0e4f26",
  1948 => x"f40e5c5b",
  1949 => x"d84c7186",
  1950 => x"ffc34a66",
  1951 => x"4ba4c29a",
  1952 => x"73496c97",
  1953 => x"517249a1",
  1954 => x"6e7e6c97",
  1955 => x"c880c148",
  1956 => x"98c758a6",
  1957 => x"7058a6cc",
  1958 => x"268ef454",
  1959 => x"264b264c",
  1960 => x"1e731e4f",
  1961 => x"dffb86f4",
  1962 => x"4bbfe087",
  1963 => x"c0e0c049",
  1964 => x"87cb0299",
  1965 => x"d1c41e73",
  1966 => x"f1fe49cc",
  1967 => x"7386c487",
  1968 => x"99c0d049",
  1969 => x"87c0c102",
  1970 => x"97d6d1c4",
  1971 => x"d1c47ebf",
  1972 => x"48bf97d7",
  1973 => x"6e58a6c8",
  1974 => x"a866c448",
  1975 => x"87e8c002",
  1976 => x"97d6d1c4",
  1977 => x"d1c449bf",
  1978 => x"481181d8",
  1979 => x"c47808e0",
  1980 => x"bf97d6d1",
  1981 => x"c1486e7e",
  1982 => x"58a6c880",
  1983 => x"a6cc98c7",
  1984 => x"d6d1c458",
  1985 => x"5066c848",
  1986 => x"494bbfe4",
  1987 => x"99c0e0c0",
  1988 => x"7387cb02",
  1989 => x"e0d1c41e",
  1990 => x"87d2fd49",
  1991 => x"497386c4",
  1992 => x"0299c0d0",
  1993 => x"c487c0c1",
  1994 => x"bf97ead1",
  1995 => x"ebd1c47e",
  1996 => x"c848bf97",
  1997 => x"486e58a6",
  1998 => x"02a866c4",
  1999 => x"c487e8c0",
  2000 => x"bf97ead1",
  2001 => x"ecd1c449",
  2002 => x"e4481181",
  2003 => x"d1c47808",
  2004 => x"7ebf97ea",
  2005 => x"80c1486e",
  2006 => x"c758a6c8",
  2007 => x"58a6cc98",
  2008 => x"48ead1c4",
  2009 => x"f85066c8",
  2010 => x"7e7087ca",
  2011 => x"f487d1f8",
  2012 => x"264b268e",
  2013 => x"d1c41e4f",
  2014 => x"d3f849cc",
  2015 => x"e0d1c487",
  2016 => x"87ccf849",
  2017 => x"49e1fac1",
  2018 => x"c287ddf7",
  2019 => x"4f2687f2",
  2020 => x"c41e731e",
  2021 => x"fa49ccd1",
  2022 => x"4a7087c1",
  2023 => x"04aab7c0",
  2024 => x"c387ccc2",
  2025 => x"c905aaf0",
  2026 => x"f8c0c287",
  2027 => x"c178c148",
  2028 => x"e0c387ed",
  2029 => x"87c905aa",
  2030 => x"48fcc0c2",
  2031 => x"dec178c1",
  2032 => x"fcc0c287",
  2033 => x"87c602bf",
  2034 => x"4ba2c0c2",
  2035 => x"4b7287c2",
  2036 => x"bff8c0c2",
  2037 => x"87e0c002",
  2038 => x"b7c44973",
  2039 => x"c2c29129",
  2040 => x"4a7381d4",
  2041 => x"92c29acf",
  2042 => x"307248c1",
  2043 => x"baff4a70",
  2044 => x"98694872",
  2045 => x"87db7970",
  2046 => x"b7c44973",
  2047 => x"c2c29129",
  2048 => x"4a7381d4",
  2049 => x"92c29acf",
  2050 => x"307248c3",
  2051 => x"69484a70",
  2052 => x"c27970b0",
  2053 => x"c048fcc0",
  2054 => x"f8c0c278",
  2055 => x"c478c048",
  2056 => x"f749ccd1",
  2057 => x"4a7087f5",
  2058 => x"03aab7c0",
  2059 => x"c087f4fd",
  2060 => x"264b2648",
  2061 => x"0000004f",
  2062 => x"00000000",
  2063 => x"00000000",
  2064 => x"724ac01e",
  2065 => x"c291c449",
  2066 => x"c081d4c2",
  2067 => x"d082c179",
  2068 => x"ee04aab7",
  2069 => x"0e4f2687",
  2070 => x"5d5c5b5e",
  2071 => x"f44d710e",
  2072 => x"4a7587e6",
  2073 => x"922ab7c4",
  2074 => x"82d4c2c2",
  2075 => x"9ccf4c75",
  2076 => x"496a94c2",
  2077 => x"c32b744b",
  2078 => x"7448c29b",
  2079 => x"ff4c7030",
  2080 => x"714874bc",
  2081 => x"f37a7098",
  2082 => x"487387f6",
  2083 => x"4c264d26",
  2084 => x"4f264b26",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"00000000",
  2088 => x"00000000",
  2089 => x"00000000",
  2090 => x"00000000",
  2091 => x"00000000",
  2092 => x"00000000",
  2093 => x"00000000",
  2094 => x"00000000",
  2095 => x"00000000",
  2096 => x"00000000",
  2097 => x"00000000",
  2098 => x"00000000",
  2099 => x"00000000",
  2100 => x"00000000",
  2101 => x"48d0ff1e",
  2102 => x"7178e1c8",
  2103 => x"08d4ff48",
  2104 => x"1e4f2678",
  2105 => x"c848d0ff",
  2106 => x"487178e1",
  2107 => x"7808d4ff",
  2108 => x"ff4866c4",
  2109 => x"267808d4",
  2110 => x"4a711e4f",
  2111 => x"1e4966c4",
  2112 => x"deff4972",
  2113 => x"48d0ff87",
  2114 => x"fc78e0c0",
  2115 => x"1e4f268e",
  2116 => x"4b711e73",
  2117 => x"1e4966c8",
  2118 => x"e0c14a73",
  2119 => x"d8ff49a2",
  2120 => x"268efc87",
  2121 => x"1e4f264b",
  2122 => x"4b711e73",
  2123 => x"fe49e2c0",
  2124 => x"4ac787e2",
  2125 => x"d4ff4813",
  2126 => x"49727808",
  2127 => x"99718ac1",
  2128 => x"ff87f105",
  2129 => x"e0c048d0",
  2130 => x"264b2678",
  2131 => x"d0ff1e4f",
  2132 => x"78c9c848",
  2133 => x"d4ff4871",
  2134 => x"4f267808",
  2135 => x"494a711e",
  2136 => x"d0ff87eb",
  2137 => x"2678c848",
  2138 => x"1e731e4f",
  2139 => x"d2c44b71",
  2140 => x"c302bfc4",
  2141 => x"87ebc287",
  2142 => x"c848d0ff",
  2143 => x"487378c9",
  2144 => x"ffb0e0c0",
  2145 => x"c47808d4",
  2146 => x"c048f8d1",
  2147 => x"0266c878",
  2148 => x"ffc387c5",
  2149 => x"c087c249",
  2150 => x"c0d2c449",
  2151 => x"0266cc59",
  2152 => x"d5c587c6",
  2153 => x"87c44ad5",
  2154 => x"4affffcf",
  2155 => x"5ac4d2c4",
  2156 => x"48c4d2c4",
  2157 => x"4b2678c1",
  2158 => x"5e0e4f26",
  2159 => x"0e5d5c5b",
  2160 => x"d2c44d71",
  2161 => x"754bbfc0",
  2162 => x"87cb029d",
  2163 => x"c291c849",
  2164 => x"714ae0c5",
  2165 => x"c287c482",
  2166 => x"c04ae0c9",
  2167 => x"7349124c",
  2168 => x"fcd1c499",
  2169 => x"b87148bf",
  2170 => x"7808d4ff",
  2171 => x"842bb7c1",
  2172 => x"04acb7c8",
  2173 => x"d1c487e7",
  2174 => x"c848bff8",
  2175 => x"fcd1c480",
  2176 => x"264d2658",
  2177 => x"264b264c",
  2178 => x"1e731e4f",
  2179 => x"4a134b71",
  2180 => x"87cb029a",
  2181 => x"e1fe4972",
  2182 => x"9a4a1387",
  2183 => x"2687f505",
  2184 => x"1e4f264b",
  2185 => x"bff8d1c4",
  2186 => x"f8d1c449",
  2187 => x"78a1c148",
  2188 => x"a9b7c0c4",
  2189 => x"ff87db03",
  2190 => x"d1c448d4",
  2191 => x"c478bffc",
  2192 => x"49bff8d1",
  2193 => x"48f8d1c4",
  2194 => x"c478a1c1",
  2195 => x"04a9b7c0",
  2196 => x"d0ff87e5",
  2197 => x"c478c848",
  2198 => x"c048c4d2",
  2199 => x"004f2678",
  2200 => x"00000000",
  2201 => x"00000000",
  2202 => x"5f000000",
  2203 => x"0000005f",
  2204 => x"00030300",
  2205 => x"00000303",
  2206 => x"147f7f14",
  2207 => x"00147f7f",
  2208 => x"6b2e2400",
  2209 => x"00123a6b",
  2210 => x"18366a4c",
  2211 => x"0032566c",
  2212 => x"594f7e30",
  2213 => x"40683a77",
  2214 => x"07040000",
  2215 => x"00000003",
  2216 => x"3e1c0000",
  2217 => x"00004163",
  2218 => x"63410000",
  2219 => x"00001c3e",
  2220 => x"1c3e2a08",
  2221 => x"082a3e1c",
  2222 => x"3e080800",
  2223 => x"0008083e",
  2224 => x"e0800000",
  2225 => x"00000060",
  2226 => x"08080800",
  2227 => x"00080808",
  2228 => x"60000000",
  2229 => x"00000060",
  2230 => x"18306040",
  2231 => x"0103060c",
  2232 => x"597f3e00",
  2233 => x"003e7f4d",
  2234 => x"7f060400",
  2235 => x"0000007f",
  2236 => x"71634200",
  2237 => x"00464f59",
  2238 => x"49632200",
  2239 => x"00367f49",
  2240 => x"13161c18",
  2241 => x"00107f7f",
  2242 => x"45672700",
  2243 => x"00397d45",
  2244 => x"4b7e3c00",
  2245 => x"00307949",
  2246 => x"71010100",
  2247 => x"00070f79",
  2248 => x"497f3600",
  2249 => x"00367f49",
  2250 => x"494f0600",
  2251 => x"001e3f69",
  2252 => x"66000000",
  2253 => x"00000066",
  2254 => x"e6800000",
  2255 => x"00000066",
  2256 => x"14080800",
  2257 => x"00222214",
  2258 => x"14141400",
  2259 => x"00141414",
  2260 => x"14222200",
  2261 => x"00080814",
  2262 => x"51030200",
  2263 => x"00060f59",
  2264 => x"5d417f3e",
  2265 => x"001e1f55",
  2266 => x"097f7e00",
  2267 => x"007e7f09",
  2268 => x"497f7f00",
  2269 => x"00367f49",
  2270 => x"633e1c00",
  2271 => x"00414141",
  2272 => x"417f7f00",
  2273 => x"001c3e63",
  2274 => x"497f7f00",
  2275 => x"00414149",
  2276 => x"097f7f00",
  2277 => x"00010109",
  2278 => x"417f3e00",
  2279 => x"007a7b49",
  2280 => x"087f7f00",
  2281 => x"007f7f08",
  2282 => x"7f410000",
  2283 => x"0000417f",
  2284 => x"40602000",
  2285 => x"003f7f40",
  2286 => x"1c087f7f",
  2287 => x"00416336",
  2288 => x"407f7f00",
  2289 => x"00404040",
  2290 => x"0c067f7f",
  2291 => x"007f7f06",
  2292 => x"0c067f7f",
  2293 => x"007f7f18",
  2294 => x"417f3e00",
  2295 => x"003e7f41",
  2296 => x"097f7f00",
  2297 => x"00060f09",
  2298 => x"61417f3e",
  2299 => x"00407e7f",
  2300 => x"097f7f00",
  2301 => x"00667f19",
  2302 => x"4d6f2600",
  2303 => x"00327b59",
  2304 => x"7f010100",
  2305 => x"0001017f",
  2306 => x"407f3f00",
  2307 => x"003f7f40",
  2308 => x"703f0f00",
  2309 => x"000f3f70",
  2310 => x"18307f7f",
  2311 => x"007f7f30",
  2312 => x"1c366341",
  2313 => x"4163361c",
  2314 => x"7c060301",
  2315 => x"0103067c",
  2316 => x"4d597161",
  2317 => x"00414347",
  2318 => x"7f7f0000",
  2319 => x"00004141",
  2320 => x"0c060301",
  2321 => x"40603018",
  2322 => x"41410000",
  2323 => x"00007f7f",
  2324 => x"03060c08",
  2325 => x"00080c06",
  2326 => x"80808080",
  2327 => x"00808080",
  2328 => x"03000000",
  2329 => x"00000407",
  2330 => x"54742000",
  2331 => x"00787c54",
  2332 => x"447f7f00",
  2333 => x"00387c44",
  2334 => x"447c3800",
  2335 => x"00004444",
  2336 => x"447c3800",
  2337 => x"007f7f44",
  2338 => x"547c3800",
  2339 => x"00185c54",
  2340 => x"7f7e0400",
  2341 => x"00000505",
  2342 => x"a4bc1800",
  2343 => x"007cfca4",
  2344 => x"047f7f00",
  2345 => x"00787c04",
  2346 => x"3d000000",
  2347 => x"0000407d",
  2348 => x"80808000",
  2349 => x"00007dfd",
  2350 => x"107f7f00",
  2351 => x"00446c38",
  2352 => x"3f000000",
  2353 => x"0000407f",
  2354 => x"180c7c7c",
  2355 => x"00787c0c",
  2356 => x"047c7c00",
  2357 => x"00787c04",
  2358 => x"447c3800",
  2359 => x"00387c44",
  2360 => x"24fcfc00",
  2361 => x"00183c24",
  2362 => x"243c1800",
  2363 => x"00fcfc24",
  2364 => x"047c7c00",
  2365 => x"00080c04",
  2366 => x"545c4800",
  2367 => x"00207454",
  2368 => x"7f3f0400",
  2369 => x"00004444",
  2370 => x"407c3c00",
  2371 => x"007c7c40",
  2372 => x"603c1c00",
  2373 => x"001c3c60",
  2374 => x"30607c3c",
  2375 => x"003c7c60",
  2376 => x"10386c44",
  2377 => x"00446c38",
  2378 => x"e0bc1c00",
  2379 => x"001c3c60",
  2380 => x"74644400",
  2381 => x"00444c5c",
  2382 => x"3e080800",
  2383 => x"00414177",
  2384 => x"7f000000",
  2385 => x"0000007f",
  2386 => x"77414100",
  2387 => x"0008083e",
  2388 => x"03010102",
  2389 => x"00010202",
  2390 => x"7f7f7f7f",
  2391 => x"007f7f7f",
  2392 => x"1c1c0808",
  2393 => x"7f7f3e3e",
  2394 => x"3e3e7f7f",
  2395 => x"08081c1c",
  2396 => x"7c181000",
  2397 => x"0010187c",
  2398 => x"7c301000",
  2399 => x"0010307c",
  2400 => x"60603010",
  2401 => x"00061e78",
  2402 => x"183c6642",
  2403 => x"0042663c",
  2404 => x"c26a3878",
  2405 => x"00386cc6",
  2406 => x"60000060",
  2407 => x"00600000",
  2408 => x"5c5b5e0e",
  2409 => x"86fc0e5d",
  2410 => x"d2c47e71",
  2411 => x"c04cbfd8",
  2412 => x"c41ec04b",
  2413 => x"c402ab66",
  2414 => x"c24dc087",
  2415 => x"754dc187",
  2416 => x"ee49731e",
  2417 => x"86c887e3",
  2418 => x"ef49e0c0",
  2419 => x"a4c487ec",
  2420 => x"f0496a4a",
  2421 => x"caf187f3",
  2422 => x"c184cc87",
  2423 => x"abb7c883",
  2424 => x"87cdff04",
  2425 => x"4d268efc",
  2426 => x"4b264c26",
  2427 => x"711e4f26",
  2428 => x"dcd2c44a",
  2429 => x"dcd2c45a",
  2430 => x"4978c748",
  2431 => x"2687e1fe",
  2432 => x"1e731e4f",
  2433 => x"b7c04a71",
  2434 => x"87d303aa",
  2435 => x"bfdce6c2",
  2436 => x"c187c405",
  2437 => x"c087c24b",
  2438 => x"e0e6c24b",
  2439 => x"c287c45b",
  2440 => x"c25ae0e6",
  2441 => x"4abfdce6",
  2442 => x"c0c19ac1",
  2443 => x"ebec49a2",
  2444 => x"c248fc87",
  2445 => x"78bfdce6",
  2446 => x"4f264b26",
  2447 => x"dce6c21e",
  2448 => x"4f2648bf",
  2449 => x"c44a711e",
  2450 => x"49721e66",
  2451 => x"fc87c0eb",
  2452 => x"1e4f268e",
  2453 => x"c348d4ff",
  2454 => x"d0ff78ff",
  2455 => x"78e1c048",
  2456 => x"c148d4ff",
  2457 => x"c4487178",
  2458 => x"08d4ff30",
  2459 => x"48d0ff78",
  2460 => x"2678e0c0",
  2461 => x"e6c21e4f",
  2462 => x"c149bfdc",
  2463 => x"c487fcd4",
  2464 => x"e848d0d2",
  2465 => x"d2c478bf",
  2466 => x"bfec48cc",
  2467 => x"d0d2c478",
  2468 => x"c3494abf",
  2469 => x"b7c899ff",
  2470 => x"7148722a",
  2471 => x"d8d2c4b0",
  2472 => x"0e4f2658",
  2473 => x"5d5c5b5e",
  2474 => x"ff4b710e",
  2475 => x"d2c487c7",
  2476 => x"50c048c8",
  2477 => x"dee64973",
  2478 => x"4c497087",
  2479 => x"eecb9cc2",
  2480 => x"87e0cb49",
  2481 => x"d2c44d70",
  2482 => x"05bf97c8",
  2483 => x"d087e2c1",
  2484 => x"d2c44966",
  2485 => x"0599bfd4",
  2486 => x"66d487d6",
  2487 => x"ccd2c449",
  2488 => x"cb0599bf",
  2489 => x"e5497387",
  2490 => x"987087ed",
  2491 => x"87c1c102",
  2492 => x"c0fe4cc1",
  2493 => x"ca497587",
  2494 => x"987087f6",
  2495 => x"c487c602",
  2496 => x"c148c8d2",
  2497 => x"c8d2c450",
  2498 => x"c005bf97",
  2499 => x"d2c487e3",
  2500 => x"d049bfd4",
  2501 => x"ff059966",
  2502 => x"d2c487d6",
  2503 => x"d449bfcc",
  2504 => x"ff059966",
  2505 => x"497387ca",
  2506 => x"7087ece4",
  2507 => x"fffe0598",
  2508 => x"26487487",
  2509 => x"264c264d",
  2510 => x"0e4f264b",
  2511 => x"5d5c5b5e",
  2512 => x"c086f80e",
  2513 => x"bfec4c4d",
  2514 => x"48a6c47e",
  2515 => x"bfd8d2c4",
  2516 => x"c01ec178",
  2517 => x"fd49c71e",
  2518 => x"86c887c9",
  2519 => x"cd029870",
  2520 => x"fa49ff87",
  2521 => x"dac187db",
  2522 => x"87ebe349",
  2523 => x"d2c44dc1",
  2524 => x"02bf97c8",
  2525 => x"e6c287cf",
  2526 => x"c149bfd4",
  2527 => x"d8e6c2b9",
  2528 => x"cefb7159",
  2529 => x"d0d2c487",
  2530 => x"e6c24bbf",
  2531 => x"c005bfdc",
  2532 => x"fdc387e9",
  2533 => x"87ffe249",
  2534 => x"e249fac3",
  2535 => x"497387f9",
  2536 => x"7199ffc3",
  2537 => x"fa49c01e",
  2538 => x"497387da",
  2539 => x"7129b7c8",
  2540 => x"fa49c11e",
  2541 => x"86c887ce",
  2542 => x"c487f4c5",
  2543 => x"4bbfd4d2",
  2544 => x"87dd029b",
  2545 => x"bfd8e6c2",
  2546 => x"87e4c749",
  2547 => x"c4059870",
  2548 => x"d24bc087",
  2549 => x"49e0c287",
  2550 => x"c287c9c7",
  2551 => x"c658dce6",
  2552 => x"d8e6c287",
  2553 => x"7378c048",
  2554 => x"0599c249",
  2555 => x"ebc387cd",
  2556 => x"87e3e149",
  2557 => x"99c24970",
  2558 => x"fb87c202",
  2559 => x"c149734c",
  2560 => x"87cd0599",
  2561 => x"e149f4c3",
  2562 => x"497087cd",
  2563 => x"c20299c2",
  2564 => x"734cfa87",
  2565 => x"0599c849",
  2566 => x"f5c387cd",
  2567 => x"87f7e049",
  2568 => x"99c24970",
  2569 => x"c487d502",
  2570 => x"02bfdcd2",
  2571 => x"c14887ca",
  2572 => x"e0d2c488",
  2573 => x"87c2c058",
  2574 => x"4dc14cff",
  2575 => x"99c44973",
  2576 => x"c387cd05",
  2577 => x"cee049f2",
  2578 => x"c2497087",
  2579 => x"87dc0299",
  2580 => x"bfdcd2c4",
  2581 => x"b7c7487e",
  2582 => x"cbc003a8",
  2583 => x"c1486e87",
  2584 => x"e0d2c480",
  2585 => x"87c2c058",
  2586 => x"4dc14cfe",
  2587 => x"ff49fdc3",
  2588 => x"7087e4df",
  2589 => x"0299c249",
  2590 => x"d2c487d5",
  2591 => x"c002bfdc",
  2592 => x"d2c487c9",
  2593 => x"78c048dc",
  2594 => x"fd87c2c0",
  2595 => x"c34dc14c",
  2596 => x"dfff49fa",
  2597 => x"497087c1",
  2598 => x"c00299c2",
  2599 => x"d2c487d9",
  2600 => x"c748bfdc",
  2601 => x"c003a8b7",
  2602 => x"d2c487c9",
  2603 => x"78c748dc",
  2604 => x"fc87c2c0",
  2605 => x"c04dc14c",
  2606 => x"c003acb7",
  2607 => x"66c487d3",
  2608 => x"80e0c148",
  2609 => x"bf6e7e70",
  2610 => x"87c5c002",
  2611 => x"7349744b",
  2612 => x"c31ec00f",
  2613 => x"dac11ef0",
  2614 => x"87c7f749",
  2615 => x"987086c8",
  2616 => x"87d8c002",
  2617 => x"bfdcd2c4",
  2618 => x"cc496e7e",
  2619 => x"4a66c491",
  2620 => x"026a8271",
  2621 => x"4b87c5c0",
  2622 => x"0f73496e",
  2623 => x"c0029d75",
  2624 => x"d2c487c8",
  2625 => x"f249bfdc",
  2626 => x"e6c287d6",
  2627 => x"c002bfe0",
  2628 => x"c24987dd",
  2629 => x"987087da",
  2630 => x"87d3c002",
  2631 => x"bfdcd2c4",
  2632 => x"87fcf149",
  2633 => x"d8f349c0",
  2634 => x"e0e6c287",
  2635 => x"f878c048",
  2636 => x"264d268e",
  2637 => x"264b264c",
  2638 => x"5b5e0e4f",
  2639 => x"fc0e5d5c",
  2640 => x"c44c7186",
  2641 => x"49bfd8d2",
  2642 => x"4da1d4c1",
  2643 => x"6981d8c1",
  2644 => x"029c747e",
  2645 => x"a5c487cf",
  2646 => x"c47b744b",
  2647 => x"49bfd8d2",
  2648 => x"6e87cbf2",
  2649 => x"059c747b",
  2650 => x"4bc087c4",
  2651 => x"4bc187c2",
  2652 => x"ccf24973",
  2653 => x"0266d487",
  2654 => x"c04987c8",
  2655 => x"4a7087e6",
  2656 => x"4ac087c2",
  2657 => x"5ae4e6c2",
  2658 => x"4d268efc",
  2659 => x"4b264c26",
  2660 => x"00004f26",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"ff4a711e",
  2666 => x"7249bfc8",
  2667 => x"4f2648a1",
  2668 => x"bfc8ff1e",
  2669 => x"c0c0fe89",
  2670 => x"a9c0c0c0",
  2671 => x"c087c401",
  2672 => x"c187c24a",
  2673 => x"2648724a",
  2674 => x"5b5e0e4f",
  2675 => x"710e5d5c",
  2676 => x"4cd4ff4b",
  2677 => x"c04866d0",
  2678 => x"ff49d678",
  2679 => x"c387f5db",
  2680 => x"496c7cff",
  2681 => x"7199ffc3",
  2682 => x"f0c3494d",
  2683 => x"a9e0c199",
  2684 => x"c387cb05",
  2685 => x"486c7cff",
  2686 => x"66d098c3",
  2687 => x"ffc37808",
  2688 => x"494a6c7c",
  2689 => x"ffc331c8",
  2690 => x"714a6c7c",
  2691 => x"c84972b2",
  2692 => x"7cffc331",
  2693 => x"b2714a6c",
  2694 => x"31c84972",
  2695 => x"6c7cffc3",
  2696 => x"ffb2714a",
  2697 => x"e0c048d0",
  2698 => x"029b7378",
  2699 => x"7b7287c2",
  2700 => x"4d264875",
  2701 => x"4b264c26",
  2702 => x"261e4f26",
  2703 => x"5b5e0e4f",
  2704 => x"86f80e5c",
  2705 => x"a6c81e76",
  2706 => x"87fdfd49",
  2707 => x"4b7086c4",
  2708 => x"a8c4486e",
  2709 => x"87f4c203",
  2710 => x"f0c34a73",
  2711 => x"aad0c19a",
  2712 => x"c187c702",
  2713 => x"c205aae0",
  2714 => x"497387e2",
  2715 => x"c30299c8",
  2716 => x"87c6ff87",
  2717 => x"9cc34c73",
  2718 => x"c105acc2",
  2719 => x"66c487c4",
  2720 => x"7131c949",
  2721 => x"4a66c41e",
  2722 => x"c492c8c1",
  2723 => x"7249e0d2",
  2724 => x"f7c3fe81",
  2725 => x"ff49d887",
  2726 => x"c887f9d8",
  2727 => x"ffc31ec0",
  2728 => x"dbfd49e0",
  2729 => x"d0ff87c1",
  2730 => x"78e0c048",
  2731 => x"1ee0ffc3",
  2732 => x"c14a66cc",
  2733 => x"d2c492c8",
  2734 => x"817249e0",
  2735 => x"87c6fffd",
  2736 => x"acc186cc",
  2737 => x"87c4c105",
  2738 => x"c94966c4",
  2739 => x"c41e7131",
  2740 => x"c8c14a66",
  2741 => x"e0d2c492",
  2742 => x"fe817249",
  2743 => x"c387edc2",
  2744 => x"c81ee0ff",
  2745 => x"c8c14a66",
  2746 => x"e0d2c492",
  2747 => x"fd817249",
  2748 => x"d787c4fd",
  2749 => x"dbd7ff49",
  2750 => x"1ec0c887",
  2751 => x"49e0ffc3",
  2752 => x"87c0d9fd",
  2753 => x"d0ff86cc",
  2754 => x"78e0c048",
  2755 => x"4c268ef8",
  2756 => x"4f264b26",
  2757 => x"5c5b5e0e",
  2758 => x"4a710e5d",
  2759 => x"d04cd4ff",
  2760 => x"b7c34d66",
  2761 => x"87c506ad",
  2762 => x"e2c148c0",
  2763 => x"751e7287",
  2764 => x"93c8c14b",
  2765 => x"83e0d2c4",
  2766 => x"f5fd4973",
  2767 => x"83c887f5",
  2768 => x"d0ff4b6b",
  2769 => x"78e1c848",
  2770 => x"48737cdd",
  2771 => x"7098ffc3",
  2772 => x"c849737c",
  2773 => x"487129b7",
  2774 => x"7098ffc3",
  2775 => x"d049737c",
  2776 => x"487129b7",
  2777 => x"7098ffc3",
  2778 => x"d848737c",
  2779 => x"7c7028b7",
  2780 => x"7c7c7cc0",
  2781 => x"7c7c7c7c",
  2782 => x"7c7c7c7c",
  2783 => x"48d0ff7c",
  2784 => x"7578e0c0",
  2785 => x"ff49dc1e",
  2786 => x"c887eed5",
  2787 => x"26487386",
  2788 => x"264c264d",
  2789 => x"1e4f264b",
  2790 => x"86fc1e73",
  2791 => x"f0c04b71",
  2792 => x"ecc04aa3",
  2793 => x"826949a3",
  2794 => x"695266cc",
  2795 => x"7080c148",
  2796 => x"98cf487e",
  2797 => x"8efc7970",
  2798 => x"4f264b26",
  2799 => x"5c5b5e0e",
  2800 => x"e94b710e",
  2801 => x"4c7087f6",
  2802 => x"87fcc6ff",
  2803 => x"c24966cc",
  2804 => x"dc0299c0",
  2805 => x"059c7487",
  2806 => x"e0c387ca",
  2807 => x"fe49731e",
  2808 => x"86c487f5",
  2809 => x"c41ee0c3",
  2810 => x"ff49ccd1",
  2811 => x"c487ffc9",
  2812 => x"4966cc86",
  2813 => x"0299c0c4",
  2814 => x"9c7487dc",
  2815 => x"c387ca05",
  2816 => x"49731ef0",
  2817 => x"c487d0fe",
  2818 => x"1ef0c386",
  2819 => x"49ccd1c4",
  2820 => x"87dac9ff",
  2821 => x"9c7486c4",
  2822 => x"cc87cf05",
  2823 => x"ffc14966",
  2824 => x"731e7199",
  2825 => x"87effd49",
  2826 => x"66cc86c4",
  2827 => x"99ffc149",
  2828 => x"d1c41e71",
  2829 => x"c8ff49cc",
  2830 => x"c5ff87f4",
  2831 => x"8efc87c2",
  2832 => x"4b264c26",
  2833 => x"5e0e4f26",
  2834 => x"fc0e5c5b",
  2835 => x"f7c4ff86",
  2836 => x"c8f3c287",
  2837 => x"d7f549bf",
  2838 => x"02987087",
  2839 => x"c487dcc1",
  2840 => x"48bfecd7",
  2841 => x"bff0d7c4",
  2842 => x"cec102a8",
  2843 => x"f4d7c487",
  2844 => x"ecd7c449",
  2845 => x"4c1181bf",
  2846 => x"aae0c34a",
  2847 => x"c387c602",
  2848 => x"c405aaf0",
  2849 => x"c24bc487",
  2850 => x"734bcf87",
  2851 => x"87d4f449",
  2852 => x"58ccf3c2",
  2853 => x"c848d0ff",
  2854 => x"d4ff78e1",
  2855 => x"7478c548",
  2856 => x"08d4ff48",
  2857 => x"48d0ff78",
  2858 => x"c478e0c0",
  2859 => x"48bfecd7",
  2860 => x"7e7080c1",
  2861 => x"c498cf48",
  2862 => x"ff58f0d7",
  2863 => x"fc87c1c3",
  2864 => x"264c268e",
  2865 => x"004f264b",
  2866 => x"00000000",
  2867 => x"5c5b5e0e",
  2868 => x"dcff0e5d",
  2869 => x"c47ec086",
  2870 => x"49bfc8d7",
  2871 => x"1e7181c2",
  2872 => x"4ac61e72",
  2873 => x"87ebd0fd",
  2874 => x"4a264871",
  2875 => x"a6cc4926",
  2876 => x"c8d7c458",
  2877 => x"81c449bf",
  2878 => x"1e721e71",
  2879 => x"d0fd4ac6",
  2880 => x"487187d1",
  2881 => x"49264a26",
  2882 => x"fc58a6d0",
  2883 => x"fec287f8",
  2884 => x"f249bfdc",
  2885 => x"987087da",
  2886 => x"87f2c902",
  2887 => x"f249e0c0",
  2888 => x"fec287c2",
  2889 => x"4cc058e0",
  2890 => x"91c44974",
  2891 => x"6981d0fe",
  2892 => x"c449744a",
  2893 => x"81bfc8d7",
  2894 => x"d7c491c4",
  2895 => x"797281d4",
  2896 => x"87d2029a",
  2897 => x"89c14972",
  2898 => x"486e9a71",
  2899 => x"7e7080c1",
  2900 => x"ff059a72",
  2901 => x"84c187ee",
  2902 => x"04acb7c2",
  2903 => x"6e87c9ff",
  2904 => x"b7fcc048",
  2905 => x"e5c804a8",
  2906 => x"744cc087",
  2907 => x"8266c84a",
  2908 => x"d7c492c4",
  2909 => x"497482d4",
  2910 => x"c48166cc",
  2911 => x"d4d7c491",
  2912 => x"694a6a81",
  2913 => x"74b97249",
  2914 => x"c8d7c44b",
  2915 => x"93c483bf",
  2916 => x"83d4d7c4",
  2917 => x"4872ba6b",
  2918 => x"a6d89871",
  2919 => x"c4497458",
  2920 => x"81bfc8d7",
  2921 => x"d7c491c4",
  2922 => x"7e6981d4",
  2923 => x"c048a6d8",
  2924 => x"5ca6d478",
  2925 => x"df4966d4",
  2926 => x"e0c60229",
  2927 => x"4a66d087",
  2928 => x"d892e0c0",
  2929 => x"ffc08266",
  2930 => x"70887248",
  2931 => x"48a6dc4a",
  2932 => x"80c478c0",
  2933 => x"4c6e78c0",
  2934 => x"d7c42cdf",
  2935 => x"78c148c4",
  2936 => x"31c34972",
  2937 => x"b1722ab7",
  2938 => x"c499ffc0",
  2939 => x"d8f0c391",
  2940 => x"6d85714d",
  2941 => x"c0c4494b",
  2942 => x"d60299c0",
  2943 => x"029c7487",
  2944 => x"c887c7c0",
  2945 => x"c578c080",
  2946 => x"d7c487d3",
  2947 => x"78c148cc",
  2948 => x"7487cac5",
  2949 => x"87d8029c",
  2950 => x"c0c24973",
  2951 => x"c00299c0",
  2952 => x"b7d087c3",
  2953 => x"fd486d2b",
  2954 => x"7098ffff",
  2955 => x"87f8c07d",
  2956 => x"bfccd7c4",
  2957 => x"87f0c002",
  2958 => x"b7d04873",
  2959 => x"58a6c828",
  2960 => x"c0029870",
  2961 => x"d7c487e2",
  2962 => x"c049bfd0",
  2963 => x"0299c0e0",
  2964 => x"7087cac0",
  2965 => x"c0e0c049",
  2966 => x"cbc00299",
  2967 => x"c2486d87",
  2968 => x"70b0c0c0",
  2969 => x"4b66c47d",
  2970 => x"c0c84973",
  2971 => x"c20299c0",
  2972 => x"d7c487c9",
  2973 => x"cc4abfd0",
  2974 => x"c0029ac0",
  2975 => x"c0c487cf",
  2976 => x"d8c0028a",
  2977 => x"c0028a87",
  2978 => x"dfc187fa",
  2979 => x"c3497387",
  2980 => x"91c299ff",
  2981 => x"81ccf0c3",
  2982 => x"dec14b11",
  2983 => x"c3497387",
  2984 => x"91c299ff",
  2985 => x"81ccf0c3",
  2986 => x"4b1181c1",
  2987 => x"c0029c74",
  2988 => x"e0c087c9",
  2989 => x"78d248a6",
  2990 => x"dc87c0c1",
  2991 => x"d2c448a6",
  2992 => x"87f7c078",
  2993 => x"ffc34973",
  2994 => x"c391c299",
  2995 => x"c181ccf0",
  2996 => x"744b1181",
  2997 => x"cac0029c",
  2998 => x"a6e0c087",
  2999 => x"78d9c148",
  3000 => x"dc87d8c0",
  3001 => x"d9c548a6",
  3002 => x"87cfc078",
  3003 => x"ffc34973",
  3004 => x"c391c299",
  3005 => x"c181ccf0",
  3006 => x"744b1181",
  3007 => x"dcc0029c",
  3008 => x"ff497387",
  3009 => x"c0fcc7b9",
  3010 => x"c4487199",
  3011 => x"98bfd0d7",
  3012 => x"58d4d7c4",
  3013 => x"c49bffc3",
  3014 => x"d4c0b3c0",
  3015 => x"c7497387",
  3016 => x"7199c0fc",
  3017 => x"d0d7c448",
  3018 => x"d7c4b0bf",
  3019 => x"ffc358d4",
  3020 => x"0266dc9b",
  3021 => x"1e87cac0",
  3022 => x"49c4d7c4",
  3023 => x"c487fdf1",
  3024 => x"c41e7386",
  3025 => x"f149c4d7",
  3026 => x"86c487f2",
  3027 => x"0266e0c0",
  3028 => x"1e87cac0",
  3029 => x"49c4d7c4",
  3030 => x"c487e1f1",
  3031 => x"4866d486",
  3032 => x"a6d830c1",
  3033 => x"c1486e58",
  3034 => x"d87e7030",
  3035 => x"80c14866",
  3036 => x"c058a6dc",
  3037 => x"04a8b7e0",
  3038 => x"d087f9f8",
  3039 => x"84c14c66",
  3040 => x"04acb7c2",
  3041 => x"c487e4f7",
  3042 => x"c848c8d7",
  3043 => x"dcff7866",
  3044 => x"264d268e",
  3045 => x"264b264c",
  3046 => x"0000004f",
  3047 => x"00000000",
  3048 => x"724ac01e",
  3049 => x"c491c449",
  3050 => x"ff81d4d7",
  3051 => x"c682c179",
  3052 => x"ee04aab7",
  3053 => x"c8d7c487",
  3054 => x"4040c048",
  3055 => x"0e4f2678",
  3056 => x"0e5c5b5e",
  3057 => x"d4ff4a71",
  3058 => x"4b66cc4c",
  3059 => x"c848d0ff",
  3060 => x"7cc278c5",
  3061 => x"8bc14973",
  3062 => x"cd029971",
  3063 => x"127c1287",
  3064 => x"c149737c",
  3065 => x"0599718b",
  3066 => x"d0ff87f3",
  3067 => x"2678c448",
  3068 => x"264b264c",
  3069 => x"4a711e4f",
  3070 => x"c848d0ff",
  3071 => x"d4ff78c5",
  3072 => x"c878c348",
  3073 => x"49721ec0",
  3074 => x"87dbc5fd",
  3075 => x"c448d0ff",
  3076 => x"268efc78",
  3077 => x"d0ff1e4f",
  3078 => x"78c5c848",
  3079 => x"c648d4ff",
  3080 => x"ff487178",
  3081 => x"ff7808d4",
  3082 => x"78c448d0",
  3083 => x"ff1e4f26",
  3084 => x"c5c848d0",
  3085 => x"48d4ff78",
  3086 => x"d0ff78ca",
  3087 => x"2678c448",
  3088 => x"5b5e0e4f",
  3089 => x"ff0e5d5c",
  3090 => x"7e7186d4",
  3091 => x"81ca496e",
  3092 => x"48496997",
  3093 => x"d428b7c5",
  3094 => x"496e58a6",
  3095 => x"699781c1",
  3096 => x"b7c54849",
  3097 => x"58a6d828",
  3098 => x"48bf976e",
  3099 => x"df58a6dc",
  3100 => x"c0c0d099",
  3101 => x"c24a6e91",
  3102 => x"c0481282",
  3103 => x"7058a6e0",
  3104 => x"92c0c44a",
  3105 => x"6e49a172",
  3106 => x"1282c34a",
  3107 => x"a6e4c048",
  3108 => x"c0807158",
  3109 => x"6e58a6e8",
  3110 => x"c880c448",
  3111 => x"66c458a6",
  3112 => x"9c4cbf97",
  3113 => x"c487c305",
  3114 => x"66d04cc0",
  3115 => x"a8b7c248",
  3116 => x"87f1cf03",
  3117 => x"c14966d0",
  3118 => x"d4c491c8",
  3119 => x"807148f0",
  3120 => x"cc58a6d0",
  3121 => x"80c84866",
  3122 => x"c858a6cc",
  3123 => x"cf02bf66",
  3124 => x"c94887d3",
  3125 => x"a6ecc028",
  3126 => x"0266d858",
  3127 => x"4d87e3c2",
  3128 => x"c3028dc3",
  3129 => x"8dc187c3",
  3130 => x"87d6c202",
  3131 => x"c4028dc4",
  3132 => x"8dc287cf",
  3133 => x"87d6c702",
  3134 => x"ca028dc8",
  3135 => x"028d87e5",
  3136 => x"cb87e6cc",
  3137 => x"87cf028d",
  3138 => x"c3028dc3",
  3139 => x"8dc287f3",
  3140 => x"87fac602",
  3141 => x"d487fccd",
  3142 => x"d3c10566",
  3143 => x"e0ffc387",
  3144 => x"c84ac04b",
  3145 => x"fefc49c0",
  3146 => x"e8c087e8",
  3147 => x"89c14966",
  3148 => x"2ad84a71",
  3149 => x"97e4ffc3",
  3150 => x"d04a715a",
  3151 => x"e5ffc32a",
  3152 => x"4a715a97",
  3153 => x"ffc32ac8",
  3154 => x"c35a97e6",
  3155 => x"5997e7ff",
  3156 => x"c280c348",
  3157 => x"f91ec450",
  3158 => x"e2f949a0",
  3159 => x"c086c487",
  3160 => x"87f1fa49",
  3161 => x"49e8d3c3",
  3162 => x"c08166d0",
  3163 => x"87f8cc51",
  3164 => x"e0fa49c2",
  3165 => x"e8d3c387",
  3166 => x"8166d049",
  3167 => x"cc51e5c0",
  3168 => x"66d487e6",
  3169 => x"c387d005",
  3170 => x"d049e8d3",
  3171 => x"51c08166",
  3172 => x"87c1fa49",
  3173 => x"c387d1cc",
  3174 => x"d049e8d3",
  3175 => x"e5c08166",
  3176 => x"f949c251",
  3177 => x"ffcb87ef",
  3178 => x"0266d487",
  3179 => x"c387cac0",
  3180 => x"d049e8d3",
  3181 => x"e5c08166",
  3182 => x"e0ffc351",
  3183 => x"c84ac04b",
  3184 => x"fcfc49c0",
  3185 => x"ffc387cc",
  3186 => x"50cb48e7",
  3187 => x"48e8d3c3",
  3188 => x"708066d0",
  3189 => x"bf976e7e",
  3190 => x"c0029949",
  3191 => x"ffc387cc",
  3192 => x"50c548e2",
  3193 => x"976e80c9",
  3194 => x"1ec950bf",
  3195 => x"49e0ffc3",
  3196 => x"c487ccf7",
  3197 => x"f849c086",
  3198 => x"486e87db",
  3199 => x"e7ca50c0",
  3200 => x"0566d487",
  3201 => x"d887f5c2",
  3202 => x"e8c04866",
  3203 => x"c0c105a8",
  3204 => x"4966dc87",
  3205 => x"c0c0c0c1",
  3206 => x"e0c091c0",
  3207 => x"c0d04a66",
  3208 => x"a17292c0",
  3209 => x"9766c449",
  3210 => x"c0c44abf",
  3211 => x"49a17292",
  3212 => x"82c54a6e",
  3213 => x"c04a6a97",
  3214 => x"7248a6e4",
  3215 => x"496e78a1",
  3216 => x"699781c7",
  3217 => x"91c0c449",
  3218 => x"82c84a6e",
  3219 => x"a14a6a97",
  3220 => x"c049744c",
  3221 => x"c08166e4",
  3222 => x"01a966e8",
  3223 => x"c087cbc1",
  3224 => x"c94966e4",
  3225 => x"d01e7131",
  3226 => x"e4fd4966",
  3227 => x"86c487de",
  3228 => x"8cc14974",
  3229 => x"c0029971",
  3230 => x"66cc87df",
  3231 => x"751ec04d",
  3232 => x"f2defd49",
  3233 => x"751ec187",
  3234 => x"caddfd49",
  3235 => x"7486c887",
  3236 => x"718cc149",
  3237 => x"e4ff0599",
  3238 => x"f549c087",
  3239 => x"d3c387f7",
  3240 => x"66d049e8",
  3241 => x"c751c081",
  3242 => x"49c287fe",
  3243 => x"c387e6f5",
  3244 => x"d049e8d3",
  3245 => x"e1c08166",
  3246 => x"87ecc751",
  3247 => x"d4f549c2",
  3248 => x"e8d3c387",
  3249 => x"8166d049",
  3250 => x"c751e5c0",
  3251 => x"66d487da",
  3252 => x"87fdc205",
  3253 => x"c04866d8",
  3254 => x"c105a8ea",
  3255 => x"66dc87c0",
  3256 => x"c0c0c149",
  3257 => x"c091c0c0",
  3258 => x"d04a66e0",
  3259 => x"7292c0c0",
  3260 => x"66c449a1",
  3261 => x"c44abf97",
  3262 => x"a17292c0",
  3263 => x"c54a6e49",
  3264 => x"4a6a9782",
  3265 => x"48a6e4c0",
  3266 => x"6e78a172",
  3267 => x"9781c749",
  3268 => x"c0c44969",
  3269 => x"c84a6e91",
  3270 => x"4a6a9782",
  3271 => x"49744ca1",
  3272 => x"8166e4c0",
  3273 => x"a966e8c0",
  3274 => x"87d3c101",
  3275 => x"c0029c74",
  3276 => x"66cc87fc",
  3277 => x"66e4c04d",
  3278 => x"7131c949",
  3279 => x"fd49751e",
  3280 => x"c387c9e1",
  3281 => x"f249e0ff",
  3282 => x"ffc387eb",
  3283 => x"49751ee0",
  3284 => x"87f2dcfd",
  3285 => x"49751ec1",
  3286 => x"87fbd9fd",
  3287 => x"e4c086cc",
  3288 => x"80c14866",
  3289 => x"58a6e8c0",
  3290 => x"ff058cc1",
  3291 => x"49c087c7",
  3292 => x"c387e2f2",
  3293 => x"d049e8d3",
  3294 => x"51c08166",
  3295 => x"c287e9c4",
  3296 => x"87d1f249",
  3297 => x"49e8d3c3",
  3298 => x"c08166d0",
  3299 => x"d7c451e1",
  3300 => x"f149c287",
  3301 => x"d3c387ff",
  3302 => x"66d049e8",
  3303 => x"51e5c081",
  3304 => x"c387c5c4",
  3305 => x"c04be0ff",
  3306 => x"49c0c84a",
  3307 => x"87e2f4fc",
  3308 => x"48e2ffc3",
  3309 => x"497450c2",
  3310 => x"ffc389c5",
  3311 => x"c35997e8",
  3312 => x"c348f4d2",
  3313 => x"2049e8ff",
  3314 => x"c3412041",
  3315 => x"c348c0d3",
  3316 => x"2049f0ff",
  3317 => x"20412041",
  3318 => x"d0412041",
  3319 => x"f0c04966",
  3320 => x"c2c0c481",
  3321 => x"d3c35997",
  3322 => x"c0c448d4",
  3323 => x"412049c0",
  3324 => x"48dcd3c3",
  3325 => x"49c4c0c4",
  3326 => x"41204120",
  3327 => x"c00266d4",
  3328 => x"ffc387c7",
  3329 => x"ffc148e0",
  3330 => x"c1497450",
  3331 => x"c31e7129",
  3332 => x"ee49e0ff",
  3333 => x"86c487e9",
  3334 => x"f8ef49c0",
  3335 => x"e8d3c387",
  3336 => x"8166d049",
  3337 => x"ffc151c0",
  3338 => x"0566d487",
  3339 => x"c387d2c1",
  3340 => x"c04be0ff",
  3341 => x"49c0c84a",
  3342 => x"87d6f2fc",
  3343 => x"48e3ffc3",
  3344 => x"e8c050c8",
  3345 => x"29d04966",
  3346 => x"97e9ffc3",
  3347 => x"66e8c059",
  3348 => x"c329c849",
  3349 => x"5997eaff",
  3350 => x"c080c148",
  3351 => x"c25066e8",
  3352 => x"49745080",
  3353 => x"1e7129c1",
  3354 => x"ed49a0f5",
  3355 => x"86c487d1",
  3356 => x"e0ee49c0",
  3357 => x"e8d3c387",
  3358 => x"8166d049",
  3359 => x"e7c051c0",
  3360 => x"e8d3c387",
  3361 => x"8166d049",
  3362 => x"c251e5c0",
  3363 => x"87c5ee49",
  3364 => x"c387d5c0",
  3365 => x"d049e8d3",
  3366 => x"e0c08166",
  3367 => x"ed49c251",
  3368 => x"c3c087f3",
  3369 => x"87c6ee87",
  3370 => x"268ed4ff",
  3371 => x"264c264d",
  3372 => x"004f264b",
  3373 => x"34364354",
  3374 => x"20202020",
  3375 => x"00000000",
  3376 => x"694d6544",
  3377 => x"66695453",
  3378 => x"44482079",
  3379 => x"20302044",
  3380 => x"00000000",
  3381 => x"20323338",
  3382 => x"00000000",
  3383 => x"32313032",
  3384 => x"39323930",
  3385 => x"00000009",
  3386 => x"731e0000",
  3387 => x"ff86e01e",
  3388 => x"c5c848d0",
  3389 => x"48d4ff78",
  3390 => x"1ed078c5",
  3391 => x"494ba6c4",
  3392 => x"87e3f1fc",
  3393 => x"d0ff86c4",
  3394 => x"ca78c448",
  3395 => x"c1496697",
  3396 => x"87c50299",
  3397 => x"e8ec4973",
  3398 => x"268ee087",
  3399 => x"1e4f264b",
  3400 => x"c44ad4ff",
  3401 => x"c448c8d8",
  3402 => x"78bff4d1",
  3403 => x"ff7affc3",
  3404 => x"78c548d0",
  3405 => x"d1c47ac4",
  3406 => x"4849bff4",
  3407 => x"7a7028d8",
  3408 => x"28d04871",
  3409 => x"48717a70",
  3410 => x"7a7028c8",
  3411 => x"bff4d1c4",
  3412 => x"48d0ff7a",
  3413 => x"4f2678c4",
  3414 => x"c44ac01e",
  3415 => x"02bffcd8",
  3416 => x"c44987ca",
  3417 => x"c148fcd8",
  3418 => x"4a1178a1",
  3419 => x"c6059a72",
  3420 => x"fcd8c487",
  3421 => x"7278c048",
  3422 => x"1e4f2648",
  3423 => x"48fcd8c4",
  3424 => x"bfd8f4c3",
  3425 => x"0e4f2678",
  3426 => x"0e5c5b5e",
  3427 => x"d0ff4a71",
  3428 => x"4bd4ff4c",
  3429 => x"d5c17cc5",
  3430 => x"7b66cc7b",
  3431 => x"7cc57cc4",
  3432 => x"c17bd3c1",
  3433 => x"c87cc47b",
  3434 => x"d4c17cc5",
  3435 => x"b749c07b",
  3436 => x"87ca06aa",
  3437 => x"81c17bc0",
  3438 => x"04a9b772",
  3439 => x"7cc487f6",
  3440 => x"d3c17cc5",
  3441 => x"c47bc07b",
  3442 => x"264c267c",
  3443 => x"1e4f264b",
  3444 => x"4b711e73",
  3445 => x"97e0f3c1",
  3446 => x"b7c249bf",
  3447 => x"f3c003a9",
  3448 => x"c41e7387",
  3449 => x"fd49dccc",
  3450 => x"c487c8cb",
  3451 => x"02987086",
  3452 => x"c487e1c0",
  3453 => x"4abfe4cc",
  3454 => x"c0c32aca",
  3455 => x"87ce028a",
  3456 => x"058ac0c1",
  3457 => x"f3c187ce",
  3458 => x"50c048e0",
  3459 => x"f3c187c6",
  3460 => x"50c148e0",
  3461 => x"4f264b26",
  3462 => x"711e731e",
  3463 => x"c6029a4a",
  3464 => x"ccddc387",
  3465 => x"c378c048",
  3466 => x"49bfc8dd",
  3467 => x"87c0ceff",
  3468 => x"c4029870",
  3469 => x"49d487cd",
  3470 => x"87e8cdff",
  3471 => x"58ccddc3",
  3472 => x"bfccddc3",
  3473 => x"87fbc005",
  3474 => x"49e0d1c4",
  3475 => x"87cbdffe",
  3476 => x"04a8b7c0",
  3477 => x"d1c487ce",
  3478 => x"defe49e0",
  3479 => x"b7c087fd",
  3480 => x"87f203a8",
  3481 => x"bfccddc3",
  3482 => x"ccddc349",
  3483 => x"78a1c148",
  3484 => x"81dcf4c3",
  3485 => x"ddc34811",
  3486 => x"ddc358d4",
  3487 => x"78c048d4",
  3488 => x"c387c0c3",
  3489 => x"02bfd4dd",
  3490 => x"c487f5c1",
  3491 => x"fe49e0d1",
  3492 => x"c087c8de",
  3493 => x"cd04a8b7",
  3494 => x"d4ddc387",
  3495 => x"88c148bf",
  3496 => x"58d8ddc3",
  3497 => x"d7c487dd",
  3498 => x"ff49bfc0",
  3499 => x"7087c1cc",
  3500 => x"cec00298",
  3501 => x"e0d1c487",
  3502 => x"d3dbfe49",
  3503 => x"ccddc387",
  3504 => x"c378c048",
  3505 => x"05bfd0dd",
  3506 => x"c387f8c1",
  3507 => x"05bfd4dd",
  3508 => x"c387f0c1",
  3509 => x"49bfccdd",
  3510 => x"48ccddc3",
  3511 => x"c378a1c1",
  3512 => x"1181dcf4",
  3513 => x"c0c2494b",
  3514 => x"ccc00299",
  3515 => x"c1487387",
  3516 => x"ddc398ff",
  3517 => x"cac158d8",
  3518 => x"d4ddc387",
  3519 => x"87c3c15b",
  3520 => x"bfd0ddc3",
  3521 => x"87fbc002",
  3522 => x"bfccddc3",
  3523 => x"ccddc349",
  3524 => x"78a1c148",
  3525 => x"81dcf4c3",
  3526 => x"1e496997",
  3527 => x"49e0d1c4",
  3528 => x"87c3dafe",
  3529 => x"ddc386c4",
  3530 => x"c148bfd0",
  3531 => x"d4ddc388",
  3532 => x"d4ddc358",
  3533 => x"c078c148",
  3534 => x"ff49ecf6",
  3535 => x"c487e5c9",
  3536 => x"2658c4d7",
  3537 => x"004f264b",
  3538 => x"00000000",
  3539 => x"00000000",
  3540 => x"00000000",
  3541 => x"00000000",
  3542 => x"711e731e",
  3543 => x"fbfd494b",
  3544 => x"d2c487e8",
  3545 => x"02bf97c8",
  3546 => x"1ec387cb",
  3547 => x"49c0c0c4",
  3548 => x"c487d4f8",
  3549 => x"fd497386",
  3550 => x"2687cffb",
  3551 => x"1e4f264b",
  3552 => x"daf61e73",
  3553 => x"49f4c787",
  3554 => x"87d8c8ff",
  3555 => x"ff494b70",
  3556 => x"7087ddc8",
  3557 => x"87cb0598",
  3558 => x"c8ff4973",
  3559 => x"987087d2",
  3560 => x"2687f502",
  3561 => x"0e4f264b",
  3562 => x"5d5c5b5e",
  3563 => x"7186f80e",
  3564 => x"fd4dc04b",
  3565 => x"7087e7d4",
  3566 => x"029b734c",
  3567 => x"c187c2c5",
  3568 => x"c148e0f3",
  3569 => x"c41e7350",
  3570 => x"fd49dccc",
  3571 => x"c487e4c3",
  3572 => x"02987086",
  3573 => x"c487ffc3",
  3574 => x"48bff4d1",
  3575 => x"d1c4b0c1",
  3576 => x"faf458f8",
  3577 => x"e0ffc387",
  3578 => x"dcccc41e",
  3579 => x"c6c9fd49",
  3580 => x"c386c487",
  3581 => x"7ebfecff",
  3582 => x"c348a6c4",
  3583 => x"78bff0ff",
  3584 => x"97e0ffc3",
  3585 => x"a9c149bf",
  3586 => x"87cac305",
  3587 => x"bfe4ffc3",
  3588 => x"71b1c149",
  3589 => x"ffcfff48",
  3590 => x"f8d1c498",
  3591 => x"e1ffc358",
  3592 => x"c248bf97",
  3593 => x"c358d8e6",
  3594 => x"49bfe8ff",
  3595 => x"87efddfd",
  3596 => x"c0029870",
  3597 => x"ffc387e2",
  3598 => x"ccc41ee0",
  3599 => x"c7fd49dc",
  3600 => x"ffc387f5",
  3601 => x"fd49bfe8",
  3602 => x"c087f4d0",
  3603 => x"f4ffc31e",
  3604 => x"87ccc449",
  3605 => x"4d7086c8",
  3606 => x"d0fd4974",
  3607 => x"1e7387e1",
  3608 => x"49dcccc4",
  3609 => x"87cbc1fd",
  3610 => x"496e86c4",
  3611 => x"87efdcfd",
  3612 => x"c0029870",
  3613 => x"ffc387e1",
  3614 => x"ccc41ee0",
  3615 => x"c6fd49dc",
  3616 => x"ffc387f5",
  3617 => x"fd49bfec",
  3618 => x"c087f4cf",
  3619 => x"c0c41ef2",
  3620 => x"cbc349c0",
  3621 => x"7486c887",
  3622 => x"e2cffd49",
  3623 => x"c41e7387",
  3624 => x"fd49dccc",
  3625 => x"c487ccc0",
  3626 => x"fd496686",
  3627 => x"7087f0db",
  3628 => x"e1c00298",
  3629 => x"e0ffc387",
  3630 => x"dcccc41e",
  3631 => x"f6c5fd49",
  3632 => x"f0ffc387",
  3633 => x"cefd49bf",
  3634 => x"f3c087f5",
  3635 => x"ccc0c41e",
  3636 => x"87ccc249",
  3637 => x"1ec286c8",
  3638 => x"49c0c0c4",
  3639 => x"c387e8f2",
  3640 => x"c0c0c41e",
  3641 => x"87dff249",
  3642 => x"d1c486c8",
  3643 => x"fe48bff4",
  3644 => x"f8d1c498",
  3645 => x"87e7f058",
  3646 => x"bfd4e6c2",
  3647 => x"d2f5fe49",
  3648 => x"f8487587",
  3649 => x"264d268e",
  3650 => x"264b264c",
  3651 => x"1e731e4f",
  3652 => x"49ca4b71",
  3653 => x"87f6dcfc",
  3654 => x"ccc41e73",
  3655 => x"fefc49dc",
  3656 => x"86c487d1",
  3657 => x"c0029870",
  3658 => x"d8c487f0",
  3659 => x"50c148c4",
  3660 => x"bfd4e6c2",
  3661 => x"c480c250",
  3662 => x"78bff4d1",
  3663 => x"50c080db",
  3664 => x"50c080cb",
  3665 => x"50c080cb",
  3666 => x"1ea0c8ff",
  3667 => x"49dcccc4",
  3668 => x"87f2c4fd",
  3669 => x"48c186c4",
  3670 => x"48c087c2",
  3671 => x"4f264b26",
  3672 => x"5c5b5e0e",
  3673 => x"86f40e5d",
  3674 => x"a6c47e71",
  3675 => x"dc78c048",
  3676 => x"f0c04d66",
  3677 => x"0266dc8d",
  3678 => x"7587e6c0",
  3679 => x"f6c1029d",
  3680 => x"8cc14c87",
  3681 => x"87efc102",
  3682 => x"d5c2028c",
  3683 => x"c2028c87",
  3684 => x"8cd087d0",
  3685 => x"87ebc402",
  3686 => x"c4028cc1",
  3687 => x"f5c487f0",
  3688 => x"c4026e87",
  3689 => x"976e87f0",
  3690 => x"e9c402bf",
  3691 => x"c41ec287",
  3692 => x"ef49c0c0",
  3693 => x"86c487d1",
  3694 => x"4bd8d8c4",
  3695 => x"49cb4a6e",
  3696 => x"87fedbfc",
  3697 => x"48e3d8c4",
  3698 => x"ccfd50c0",
  3699 => x"d8c487d0",
  3700 => x"d1c458d0",
  3701 => x"c148bff4",
  3702 => x"f8d1c4b0",
  3703 => x"87ffec58",
  3704 => x"49d8d8c4",
  3705 => x"c487e8ef",
  3706 => x"fd49d8d8",
  3707 => x"c487d6e0",
  3708 => x"78c148a6",
  3709 => x"7587dfc3",
  3710 => x"ff49c01e",
  3711 => x"7587d5c4",
  3712 => x"87fbf549",
  3713 => x"66c81e75",
  3714 => x"c7c4ff49",
  3715 => x"7586c887",
  3716 => x"91c8c149",
  3717 => x"81e0d2c4",
  3718 => x"a6c481c8",
  3719 => x"c2786948",
  3720 => x"497587f4",
  3721 => x"c491c8c1",
  3722 => x"7148e0d2",
  3723 => x"58a6c880",
  3724 => x"c84866c4",
  3725 => x"58a6cc80",
  3726 => x"c04866c8",
  3727 => x"c0026e78",
  3728 => x"4c7587e5",
  3729 => x"d8c494cc",
  3730 => x"4b7484cc",
  3731 => x"49cb4a6e",
  3732 => x"87eed9fc",
  3733 => x"c049a4cb",
  3734 => x"c81e7451",
  3735 => x"f9fc4966",
  3736 => x"86c487d1",
  3737 => x"7587cac0",
  3738 => x"c491cc49",
  3739 => x"c081ccd8",
  3740 => x"e9c9fd51",
  3741 => x"754a7087",
  3742 => x"c491c449",
  3743 => x"7281c8d8",
  3744 => x"bf66c879",
  3745 => x"87d9c002",
  3746 => x"89c24975",
  3747 => x"7148c0d0",
  3748 => x"c4497030",
  3749 => x"48bff4d1",
  3750 => x"d1c4b071",
  3751 => x"d8c058f8",
  3752 => x"c2497587",
  3753 => x"48c0d089",
  3754 => x"49703071",
  3755 => x"d1c4b9ff",
  3756 => x"7148bff4",
  3757 => x"f8d1c498",
  3758 => x"48a6c458",
  3759 => x"78bf66c8",
  3760 => x"6e87d3c0",
  3761 => x"87dff349",
  3762 => x"c058a6c8",
  3763 => x"496e87c8",
  3764 => x"c887faf8",
  3765 => x"d1c458a6",
  3766 => x"fe48bff4",
  3767 => x"f8d1c498",
  3768 => x"87fbe858",
  3769 => x"f44866c4",
  3770 => x"264d268e",
  3771 => x"264b264c",
  3772 => x"1e731e4f",
  3773 => x"48f4d1c4",
  3774 => x"f3c178c1",
  3775 => x"50c148e0",
  3776 => x"48c4c8c1",
  3777 => x"d6e850c0",
  3778 => x"c41ec387",
  3779 => x"e949c0c0",
  3780 => x"1ec287f5",
  3781 => x"49c0c0c4",
  3782 => x"c887ece9",
  3783 => x"f0f4c386",
  3784 => x"c2f249bf",
  3785 => x"05987087",
  3786 => x"e787efc1",
  3787 => x"f4c387f1",
  3788 => x"ea49bfec",
  3789 => x"f4c387d9",
  3790 => x"fd49bfec",
  3791 => x"c487c6db",
  3792 => x"48bff4d1",
  3793 => x"d1c498fe",
  3794 => x"d2e758f8",
  3795 => x"49d0c687",
  3796 => x"87d0f9fe",
  3797 => x"fe494b70",
  3798 => x"7087d5f9",
  3799 => x"87cc0598",
  3800 => x"f9fe4973",
  3801 => x"987087ca",
  3802 => x"87f4ff02",
  3803 => x"bff4d1c4",
  3804 => x"c4b0c148",
  3805 => x"e658f8d1",
  3806 => x"e4c187e5",
  3807 => x"e3f8fe49",
  3808 => x"494b7087",
  3809 => x"87e8f8fe",
  3810 => x"c0059870",
  3811 => x"497387cc",
  3812 => x"87dcf8fe",
  3813 => x"ff029870",
  3814 => x"d1c487f4",
  3815 => x"fe48bff4",
  3816 => x"f8d1c498",
  3817 => x"87f7e558",
  3818 => x"87f4cfff",
  3819 => x"87d0c7fe",
  3820 => x"e3e949c1",
  3821 => x"2648c087",
  3822 => x"1e4f264b",
  3823 => x"4b711e73",
  3824 => x"87c8c4ff",
  3825 => x"cffe4973",
  3826 => x"4b2687c6",
  3827 => x"5e0e4f26",
  3828 => x"fc0e5c5b",
  3829 => x"ffffc186",
  3830 => x"c04b6e4c",
  3831 => x"87f8e849",
  3832 => x"87d7edfe",
  3833 => x"87d5f9fe",
  3834 => x"7387ffe3",
  3835 => x"c1997449",
  3836 => x"05997183",
  3837 => x"fffd87e5",
  3838 => x"497087ea",
  3839 => x"87e7d4fe",
  3840 => x"fc87d8ff",
  3841 => x"264c268e",
  3842 => x"004f264b",
  3843 => x"f5f2ebf4",
  3844 => x"0c040605",
  3845 => x"0a830b03",
  3846 => x"00000066",
  3847 => x"00da005a",
  3848 => x"08948000",
  3849 => x"00788005",
  3850 => x"00018002",
  3851 => x"00098003",
  3852 => x"00008004",
  3853 => x"08918001",
  3854 => x"00000026",
  3855 => x"0000001d",
  3856 => x"0000001c",
  3857 => x"00000025",
  3858 => x"0000001a",
  3859 => x"0000001b",
  3860 => x"00000024",
  3861 => x"00000112",
  3862 => x"0000002e",
  3863 => x"0000002d",
  3864 => x"00000023",
  3865 => x"00000036",
  3866 => x"00000021",
  3867 => x"0000002b",
  3868 => x"0000002c",
  3869 => x"00000022",
  3870 => x"006c003d",
  3871 => x"00000035",
  3872 => x"00000034",
  3873 => x"0075003e",
  3874 => x"00000032",
  3875 => x"00000033",
  3876 => x"006b003c",
  3877 => x"0000002a",
  3878 => x"007d0046",
  3879 => x"00730043",
  3880 => x"0069003b",
  3881 => x"00ca0045",
  3882 => x"0070003a",
  3883 => x"00720042",
  3884 => x"00740044",
  3885 => x"00000031",
  3886 => x"00000055",
  3887 => x"007c004d",
  3888 => x"007a004b",
  3889 => x"0000007b",
  3890 => x"00710049",
  3891 => x"0084004c",
  3892 => x"00770054",
  3893 => x"00000041",
  3894 => x"00000061",
  3895 => x"007c005b",
  3896 => x"00000052",
  3897 => x"000000f1",
  3898 => x"00000259",
  3899 => x"005d000e",
  3900 => x"0000005d",
  3901 => x"0079004a",
  3902 => x"00000016",
  3903 => x"00070076",
  3904 => x"000d0414",
  3905 => x"0000001e",
  3906 => x"00000029",
  3907 => x"00000011",
  3908 => x"00000015",
  3909 => x"00004000",
  3910 => x"00003d34",
  3911 => x"0882ff01",
  3912 => x"64f3c8f3",
  3913 => x"01f250f3",
  3914 => x"00f40181",
  3915 => x"00003fa0",
  3916 => x"00003fac",
  3917 => x"72617441",
  3918 => x"54532069",
  3919 => x"31503b3b",
  3920 => x"6f74532c",
  3921 => x"65676172",
  3922 => x"5331503b",
  3923 => x"532c5530",
  3924 => x"462c2054",
  3925 => x"70706f6c",
  3926 => x"3a412079",
  3927 => x"5331503b",
  3928 => x"532c5531",
  3929 => x"462c2054",
  3930 => x"70706f6c",
  3931 => x"3a422079",
  3932 => x"4f31503b",
  3933 => x"572c3736",
  3934 => x"65746972",
  3935 => x"6f727020",
  3936 => x"74636574",
  3937 => x"66664f2c",
  3938 => x"2c3a412c",
  3939 => x"422c3a42",
  3940 => x"3b68746f",
  3941 => x"414f3150",
  3942 => x"61482c42",
  3943 => x"64206472",
  3944 => x"736b7369",
  3945 => x"6e6f4e2c",
  3946 => x"6e552c65",
  3947 => x"30207469",
  3948 => x"696e552c",
  3949 => x"2c312074",
  3950 => x"68746f42",
  3951 => x"5331503b",
  3952 => x"482c5532",
  3953 => x"48564644",
  3954 => x"61482c44",
  3955 => x"69666472",
  3956 => x"3020656c",
  3957 => x"5331503b",
  3958 => x"482c5533",
  3959 => x"48564644",
  3960 => x"61482c44",
  3961 => x"69666472",
  3962 => x"3120656c",
  3963 => x"2c32503b",
  3964 => x"74737953",
  3965 => x"503b6d65",
  3966 => x"4f4e4f32",
  3967 => x"6968432c",
  3968 => x"74657370",
  3969 => x"2c54532c",
  3970 => x"2c455453",
  3971 => x"6167654d",
  3972 => x"2c455453",
  3973 => x"72455453",
  3974 => x"7364696f",
  3975 => x"4f32503b",
  3976 => x"54532c4a",
  3977 => x"696c4220",
  3978 => x"72657474",
  3979 => x"66664f2c",
  3980 => x"3b6e4f2c",
  3981 => x"314f3250",
  3982 => x"41522c33",
  3983 => x"6e28204d",
  3984 => x"20646565",
  3985 => x"64726148",
  3986 => x"73655220",
  3987 => x"2c297465",
  3988 => x"4b323135",
  3989 => x"424d312c",
  3990 => x"424d322c",
  3991 => x"424d342c",
  3992 => x"424d382c",
  3993 => x"4d34312c",
  3994 => x"32503b42",
  3995 => x"4d492c46",
  3996 => x"4d4f5247",
  3997 => x"616f4c2c",
  3998 => x"4f522064",
  3999 => x"32503b4d",
  4000 => x"49422c46",
  4001 => x"4354534e",
  4002 => x"616f4c2c",
  4003 => x"61432064",
  4004 => x"69727472",
  4005 => x"3b656764",
  4006 => x"532c3350",
  4007 => x"646e756f",
  4008 => x"56202620",
  4009 => x"6f656469",
  4010 => x"4f33503b",
  4011 => x"69562c38",
  4012 => x"206f6564",
  4013 => x"65646f6d",
  4014 => x"6e6f4d2c",
  4015 => x"6f432c6f",
  4016 => x"72756f6c",
  4017 => x"4f33503b",
  4018 => x"69562c53",
  4019 => x"676e696b",
  4020 => x"314d532f",
  4021 => x"4f2c3439",
  4022 => x"4f2c6666",
  4023 => x"33503b6e",
  4024 => x"2c4c4b4f",
  4025 => x"6e616353",
  4026 => x"656e696c",
  4027 => x"664f2c73",
  4028 => x"35322c66",
  4029 => x"30352c25",
  4030 => x"35372c25",
  4031 => x"33503b25",
  4032 => x"432c544f",
  4033 => x"6f706d6f",
  4034 => x"65746973",
  4035 => x"656c6220",
  4036 => x"4f2c646e",
  4037 => x"4f2c6666",
  4038 => x"33503b6e",
  4039 => x"532c4d4f",
  4040 => x"65726574",
  4041 => x"6f73206f",
  4042 => x"2c646e75",
  4043 => x"2c66664f",
  4044 => x"503b6e4f",
  4045 => x"2c554f33",
  4046 => x"69657453",
  4047 => x"7265626e",
  4048 => x"6f642067",
  4049 => x"656c676e",
  4050 => x"66664f2c",
  4051 => x"3b6e4f2c",
  4052 => x"432c4353",
  4053 => x"4c2c4746",
  4054 => x"2064616f",
  4055 => x"666e6f63",
  4056 => x"533b6769",
  4057 => x"46432c44",
  4058 => x"61532c47",
  4059 => x"63206576",
  4060 => x"69666e6f",
  4061 => x"30543b67",
  4062 => x"7365522c",
  4063 => x"28207465",
  4064 => x"646c6f48",
  4065 => x"726f6620",
  4066 => x"72616820",
  4067 => x"65722064",
  4068 => x"29746573",
  4069 => x"762c563b",
  4070 => x"30342e33",
  4071 => x"0000002e",
  4072 => x"20534f54",
  4073 => x"20202020",
  4074 => x"00474d49",
  4075 => x"5453494d",
  4076 => x"20595245",
  4077 => x"00474643",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
